magic
tech sky130A
magscale 1 2
timestamp 1714065493
<< error_s >>
rect 3042 -1758 3808 -316
<< dnwell >>
rect 2668 -1758 3808 -316
<< locali >>
rect 2726 -315 3744 -284
rect 2726 -349 2750 -315
rect 2784 -349 2822 -315
rect 2856 -349 2894 -315
rect 2928 -349 2966 -315
rect 3000 -349 3038 -315
rect 3072 -349 3110 -315
rect 3144 -349 3182 -315
rect 3216 -349 3254 -315
rect 3288 -349 3326 -315
rect 3360 -349 3398 -315
rect 3432 -349 3470 -315
rect 3504 -349 3542 -315
rect 3576 -349 3614 -315
rect 3648 -349 3686 -315
rect 3720 -349 3744 -315
rect 2726 -380 3744 -349
rect 4622 -423 5296 -416
rect 784 -512 836 -478
rect 870 -512 908 -478
rect 942 -512 980 -478
rect 1014 -512 1052 -478
rect 1086 -512 1124 -478
rect 1158 -512 1196 -478
rect 1230 -512 1282 -478
rect 750 -574 784 -512
rect 1282 -574 1316 -512
rect 4622 -529 4654 -423
rect 5264 -529 5296 -423
rect 4622 -536 5296 -529
rect 2726 -1023 3744 -992
rect 2726 -1057 2750 -1023
rect 2784 -1057 2822 -1023
rect 2856 -1057 2894 -1023
rect 2928 -1057 2966 -1023
rect 3000 -1057 3038 -1023
rect 3072 -1057 3110 -1023
rect 3144 -1057 3182 -1023
rect 3216 -1057 3254 -1023
rect 3288 -1057 3326 -1023
rect 3360 -1057 3398 -1023
rect 3432 -1057 3470 -1023
rect 3504 -1057 3542 -1023
rect 3576 -1057 3614 -1023
rect 3648 -1057 3686 -1023
rect 3720 -1057 3744 -1023
rect 2726 -1088 3744 -1057
rect 758 -1564 792 -1502
rect 1272 -1564 1306 -1502
rect 792 -1598 835 -1564
rect 869 -1598 907 -1564
rect 941 -1598 979 -1564
rect 1013 -1598 1051 -1564
rect 1085 -1598 1123 -1564
rect 1157 -1598 1195 -1564
rect 1229 -1598 1272 -1564
rect 3984 -1551 4658 -1544
rect 3984 -1657 4016 -1551
rect 4626 -1657 4658 -1551
rect 3984 -1664 4658 -1657
rect 2728 -1729 3746 -1698
rect 2728 -1763 2752 -1729
rect 2786 -1763 2824 -1729
rect 2858 -1763 2896 -1729
rect 2930 -1763 2968 -1729
rect 3002 -1763 3040 -1729
rect 3074 -1763 3112 -1729
rect 3146 -1763 3184 -1729
rect 3218 -1763 3256 -1729
rect 3290 -1763 3328 -1729
rect 3362 -1763 3400 -1729
rect 3434 -1763 3472 -1729
rect 3506 -1763 3544 -1729
rect 3578 -1763 3616 -1729
rect 3650 -1763 3688 -1729
rect 3722 -1763 3746 -1729
rect 2728 -1794 3746 -1763
<< viali >>
rect 2750 -349 2784 -315
rect 2822 -349 2856 -315
rect 2894 -349 2928 -315
rect 2966 -349 3000 -315
rect 3038 -349 3072 -315
rect 3110 -349 3144 -315
rect 3182 -349 3216 -315
rect 3254 -349 3288 -315
rect 3326 -349 3360 -315
rect 3398 -349 3432 -315
rect 3470 -349 3504 -315
rect 3542 -349 3576 -315
rect 3614 -349 3648 -315
rect 3686 -349 3720 -315
rect 750 -512 784 -478
rect 836 -512 870 -478
rect 908 -512 942 -478
rect 980 -512 1014 -478
rect 1052 -512 1086 -478
rect 1124 -512 1158 -478
rect 1196 -512 1230 -478
rect 1282 -512 1316 -478
rect 4654 -529 5264 -423
rect 2750 -1057 2784 -1023
rect 2822 -1057 2856 -1023
rect 2894 -1057 2928 -1023
rect 2966 -1057 3000 -1023
rect 3038 -1057 3072 -1023
rect 3110 -1057 3144 -1023
rect 3182 -1057 3216 -1023
rect 3254 -1057 3288 -1023
rect 3326 -1057 3360 -1023
rect 3398 -1057 3432 -1023
rect 3470 -1057 3504 -1023
rect 3542 -1057 3576 -1023
rect 3614 -1057 3648 -1023
rect 3686 -1057 3720 -1023
rect 758 -1598 792 -1564
rect 835 -1598 869 -1564
rect 907 -1598 941 -1564
rect 979 -1598 1013 -1564
rect 1051 -1598 1085 -1564
rect 1123 -1598 1157 -1564
rect 1195 -1598 1229 -1564
rect 1272 -1598 1306 -1564
rect 4016 -1657 4626 -1551
rect 2752 -1763 2786 -1729
rect 2824 -1763 2858 -1729
rect 2896 -1763 2930 -1729
rect 2968 -1763 3002 -1729
rect 3040 -1763 3074 -1729
rect 3112 -1763 3146 -1729
rect 3184 -1763 3218 -1729
rect 3256 -1763 3290 -1729
rect 3328 -1763 3362 -1729
rect 3400 -1763 3434 -1729
rect 3472 -1763 3506 -1729
rect 3544 -1763 3578 -1729
rect 3616 -1763 3650 -1729
rect 3688 -1763 3722 -1729
<< metal1 >>
rect 652 -478 1434 -128
rect 652 -512 750 -478
rect 784 -512 836 -478
rect 870 -512 908 -478
rect 942 -512 980 -478
rect 1014 -512 1052 -478
rect 1086 -512 1124 -478
rect 1158 -512 1196 -478
rect 1230 -512 1282 -478
rect 1316 -512 1434 -478
rect 652 -526 1434 -512
rect 652 -580 796 -526
rect 960 -586 1106 -526
rect 1270 -580 1434 -526
rect 2580 -315 3852 -128
rect 2580 -349 2750 -315
rect 2784 -349 2822 -315
rect 2856 -349 2894 -315
rect 2928 -349 2966 -315
rect 3000 -349 3038 -315
rect 3072 -349 3110 -315
rect 3144 -349 3182 -315
rect 3216 -349 3254 -315
rect 3288 -349 3326 -315
rect 3360 -349 3398 -315
rect 3432 -349 3470 -315
rect 3504 -349 3542 -315
rect 3576 -349 3614 -315
rect 3648 -349 3686 -315
rect 3720 -349 3852 -315
rect 2580 -422 3852 -349
rect 932 -626 1134 -586
rect 820 -712 1472 -688
rect 820 -764 1200 -712
rect 1252 -764 1264 -712
rect 1316 -764 1328 -712
rect 1380 -764 1392 -712
rect 1444 -764 1472 -712
rect 820 -788 1472 -764
rect 820 -972 900 -788
rect 652 -1288 900 -972
rect 982 -988 1082 -850
rect 2580 -948 2772 -422
rect 2838 -499 2904 -492
rect 2838 -551 2845 -499
rect 2897 -551 2904 -499
rect 3136 -502 3336 -422
rect 3568 -499 3634 -492
rect 2838 -558 2904 -551
rect 2936 -552 3536 -502
rect 3568 -551 3575 -499
rect 3627 -551 3634 -499
rect 2846 -812 2904 -558
rect 3568 -558 3634 -551
rect 2936 -596 3534 -586
rect 2936 -776 2953 -596
rect 3517 -776 3534 -596
rect 2936 -788 3534 -776
rect 3568 -812 3626 -558
rect 2936 -868 3536 -822
rect 3136 -948 3336 -868
rect 3700 -948 3852 -422
rect 982 -1012 1472 -988
rect 982 -1064 1191 -1012
rect 1243 -1064 1255 -1012
rect 1307 -1064 1319 -1012
rect 1371 -1064 1383 -1012
rect 1435 -1064 1472 -1012
rect 982 -1088 1472 -1064
rect 2580 -1023 3852 -948
rect 2580 -1057 2750 -1023
rect 2784 -1057 2822 -1023
rect 2856 -1057 2894 -1023
rect 2928 -1057 2966 -1023
rect 3000 -1057 3038 -1023
rect 3072 -1057 3110 -1023
rect 3144 -1057 3182 -1023
rect 3216 -1057 3254 -1023
rect 3288 -1057 3326 -1023
rect 3360 -1057 3398 -1023
rect 3432 -1057 3470 -1023
rect 3504 -1057 3542 -1023
rect 3576 -1057 3614 -1023
rect 3648 -1057 3686 -1023
rect 3720 -1057 3852 -1023
rect 982 -1226 1082 -1088
rect 2580 -1132 3852 -1057
rect 652 -1356 1210 -1288
rect 820 -1388 1210 -1356
rect 932 -1492 1132 -1448
rect 652 -1552 804 -1496
rect 958 -1552 1104 -1492
rect 1260 -1552 1418 -1496
rect 652 -1564 1418 -1552
rect 652 -1598 758 -1564
rect 792 -1598 835 -1564
rect 869 -1598 907 -1564
rect 941 -1598 979 -1564
rect 1013 -1598 1051 -1564
rect 1085 -1598 1123 -1564
rect 1157 -1598 1195 -1564
rect 1229 -1598 1272 -1564
rect 1306 -1598 1418 -1564
rect 652 -1950 1418 -1598
rect 2580 -1658 2772 -1132
rect 3136 -1212 3336 -1132
rect 2936 -1258 3536 -1212
rect 2846 -1522 2904 -1268
rect 2936 -1302 3534 -1292
rect 2936 -1482 2953 -1302
rect 3517 -1482 3534 -1302
rect 2936 -1494 3534 -1482
rect 2838 -1529 2904 -1522
rect 3568 -1522 3626 -1268
rect 2838 -1581 2845 -1529
rect 2897 -1581 2904 -1529
rect 2936 -1578 3536 -1526
rect 3568 -1529 3634 -1522
rect 2838 -1588 2904 -1581
rect 3136 -1658 3336 -1578
rect 3568 -1581 3575 -1529
rect 3627 -1581 3634 -1529
rect 3568 -1588 3634 -1581
rect 3700 -1658 3852 -1132
rect 2580 -1729 3852 -1658
rect 2580 -1763 2752 -1729
rect 2786 -1763 2824 -1729
rect 2858 -1763 2896 -1729
rect 2930 -1763 2968 -1729
rect 3002 -1763 3040 -1729
rect 3074 -1763 3112 -1729
rect 3146 -1763 3184 -1729
rect 3218 -1763 3256 -1729
rect 3290 -1763 3328 -1729
rect 3362 -1763 3400 -1729
rect 3434 -1763 3472 -1729
rect 3506 -1763 3544 -1729
rect 3578 -1763 3616 -1729
rect 3650 -1763 3688 -1729
rect 3722 -1763 3852 -1729
rect 2580 -1950 3852 -1763
rect 3912 -378 5370 -128
rect 3912 -1520 4086 -378
rect 4588 -423 5370 -378
rect 4230 -448 4450 -438
rect 4230 -628 4250 -448
rect 4430 -628 4450 -448
rect 4230 -638 4450 -628
rect 4588 -529 4654 -423
rect 5264 -529 5370 -423
rect 4588 -560 5370 -529
rect 4148 -854 4528 -786
rect 4148 -1226 4248 -854
rect 4428 -1226 4528 -854
rect 4148 -1286 4528 -1226
rect 4238 -1520 4440 -1446
rect 4588 -1520 4696 -560
rect 4842 -634 5044 -560
rect 4756 -852 5136 -788
rect 4756 -1224 4852 -852
rect 5032 -1224 5136 -852
rect 4756 -1288 5136 -1224
rect 3912 -1551 4696 -1520
rect 3912 -1657 4016 -1551
rect 4626 -1657 4696 -1551
rect 4832 -1450 5052 -1440
rect 4832 -1630 4852 -1450
rect 5032 -1630 5052 -1450
rect 4832 -1640 5052 -1630
rect 3912 -1700 4696 -1657
rect 5196 -1700 5370 -560
rect 3912 -1950 5370 -1700
<< via1 >>
rect 1200 -764 1252 -712
rect 1264 -764 1316 -712
rect 1328 -764 1380 -712
rect 1392 -764 1444 -712
rect 2845 -551 2897 -499
rect 3575 -551 3627 -499
rect 2953 -776 3517 -596
rect 1191 -1064 1243 -1012
rect 1255 -1064 1307 -1012
rect 1319 -1064 1371 -1012
rect 1383 -1064 1435 -1012
rect 2953 -1482 3517 -1302
rect 2845 -1581 2897 -1529
rect 3575 -1581 3627 -1529
rect 4250 -628 4430 -448
rect 4248 -1226 4428 -854
rect 4852 -1224 5032 -852
rect 4852 -1630 5032 -1450
<< metal2 >>
rect 3742 -448 5670 -438
rect 1854 -499 3634 -452
rect 1854 -551 2845 -499
rect 2897 -551 3575 -499
rect 3627 -551 3634 -499
rect 1854 -558 3634 -551
rect 1854 -688 1954 -558
rect 1166 -712 1954 -688
rect 1166 -764 1200 -712
rect 1252 -764 1264 -712
rect 1316 -764 1328 -712
rect 1380 -764 1392 -712
rect 1444 -764 1954 -712
rect 1166 -788 1954 -764
rect 2936 -588 3534 -586
rect 3742 -588 4250 -448
rect 2936 -596 4250 -588
rect 2936 -776 2953 -596
rect 3517 -628 4250 -596
rect 4430 -628 5670 -448
rect 3517 -638 5670 -628
rect 3517 -776 3942 -638
rect 2936 -788 3942 -776
rect 4240 -854 4438 -840
rect 1152 -1012 2074 -988
rect 1152 -1064 1191 -1012
rect 1243 -1064 1255 -1012
rect 1307 -1064 1319 -1012
rect 1371 -1064 1383 -1012
rect 1435 -1064 2074 -1012
rect 1152 -1088 2074 -1064
rect 1822 -1522 2074 -1088
rect 4240 -1226 4248 -854
rect 4428 -1226 4438 -854
rect 2936 -1302 3942 -1292
rect 2936 -1482 2953 -1302
rect 3517 -1440 3942 -1302
rect 4240 -1440 4438 -1226
rect 4844 -852 5042 -638
rect 4844 -1224 4852 -852
rect 5032 -1224 5042 -852
rect 4844 -1238 5042 -1224
rect 3517 -1450 5670 -1440
rect 3517 -1482 4852 -1450
rect 2936 -1492 4852 -1482
rect 2936 -1494 3534 -1492
rect 1822 -1529 3634 -1522
rect 1822 -1581 2845 -1529
rect 2897 -1581 3575 -1529
rect 3627 -1581 3634 -1529
rect 1822 -1628 3634 -1581
rect 3742 -1630 4852 -1492
rect 5032 -1630 5670 -1450
rect 3742 -1640 5670 -1630
use sky130_fd_pr__nfet_01v8_69TQ3K  XM1 ../../chipalooza/sky130_od_ip__tempsensor/mag
timestamp 1713225924
transform 0 -1 1032 1 0 -1338
box -286 -300 286 300
use sky130_fd_pr__pfet_01v8_3HMWVM  XM2 ../../chipalooza/sky130_od_ip__tempsensor/mag
timestamp 1713225924
transform 0 -1 1033 1 0 -738
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM3
timestamp 1713225924
transform 0 1 3236 -1 0 -687
box -347 -548 347 548
use sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B  XM4
timestamp 1713225924
transform 0 1 3236 -1 0 -1393
box -347 -548 347 548
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM5
timestamp 1713225924
transform 0 1 4339 -1 0 -1040
box -658 -397 658 397
use sky130_fd_pr__pfet_g5v0d10v5_VHBZVD  XM6
timestamp 1713225924
transform 0 1 4943 -1 0 -1040
box -658 -397 658 397
<< labels >>
flabel metal1 s 652 -478 1434 -128 0 FreeSans 2000 0 0 0 dvdd
port 1 nsew
flabel metal1 s 652 -1950 1418 -1598 0 FreeSans 2000 0 0 0 dvss
port 2 nsew
flabel metal1 s 3912 -378 5370 -128 0 FreeSans 2000 0 0 0 avdd
port 3 nsew
flabel metal1 s 2580 -1950 3852 -1794 0 FreeSans 1500 0 0 0 avss
port 4 nsew
flabel metal1 s 652 -1356 900 -972 0 FreeSans 1500 0 0 0 in
port 5 nsew
flabel metal2 s 1822 -1628 2074 -988 0 FreeSans 1000 0 0 0 in_b
port 6 nsew
flabel metal2 s 4440 -638 5670 -438 0 FreeSans 1500 0 0 0 out_b
port 7 nsew
flabel metal2 s 5042 -1640 5670 -1440 0 FreeSans 1500 0 0 0 out
port 8 nsew
<< properties >>
string GDS_END 2855258
string GDS_FILE ../../chipalooza/sky130_be_ip__lsxo/gds/sky130_be_ip__lsxo.gds
string GDS_START 2834554
<< end >>
