magic
tech sky130A
magscale 1 2
timestamp 1713983242
<< dnwell >>
rect 410 30 3346 1630
rect 410 -2800 4354 30
<< nwell >>
rect 301 1424 3546 1830
rect 301 482 616 1424
rect 3204 482 3546 1424
rect 301 373 3546 482
rect 301 -2594 616 373
rect 1957 230 3546 373
rect 1957 -297 4463 230
rect 3362 -482 4463 -297
rect 4148 -2594 4463 -482
rect 301 -2911 4463 -2594
<< mvnsubdiff >>
rect 367 1744 3480 1764
rect 367 1710 447 1744
rect 3440 1710 3480 1744
rect 367 1690 3480 1710
rect 367 1684 441 1690
rect 367 -2763 387 1684
rect 421 -2763 441 1684
rect 3406 1672 3480 1690
rect 3406 200 3426 1672
rect 3460 200 3480 1672
rect 3406 164 3480 200
rect 3406 144 4397 164
rect 3406 110 3482 144
rect 4317 110 4397 144
rect 3406 90 4397 110
rect 367 -2769 441 -2763
rect 4323 84 4397 90
rect 4323 -2763 4343 84
rect 4377 -2763 4397 84
rect 4323 -2769 4397 -2763
rect 367 -2789 4397 -2769
rect 367 -2823 447 -2789
rect 4317 -2823 4397 -2789
rect 367 -2843 4397 -2823
<< mvnsubdiffcont >>
rect 447 1710 3440 1744
rect 387 -2763 421 1684
rect 3426 200 3460 1672
rect 3482 110 4317 144
rect 4343 -2763 4377 84
rect 447 -2823 4317 -2789
<< locali >>
rect 387 1710 447 1744
rect 3440 1710 3460 1744
rect 387 1684 3460 1710
rect 421 1672 3460 1684
rect 421 1621 3426 1672
rect 421 482 571 1621
rect 616 556 768 1376
rect 1169 1355 1343 1377
rect 1169 674 1221 1355
rect 1297 674 1343 1355
rect 1169 556 1343 674
rect 1753 1373 1903 1377
rect 2850 1375 3087 1376
rect 2423 1373 3087 1375
rect 1753 1357 3087 1373
rect 1753 676 1802 1357
rect 1878 1352 3087 1357
rect 1878 847 2225 1352
rect 1878 676 1927 847
rect 1753 556 1927 676
rect 2164 623 2225 847
rect 2355 1339 3087 1352
rect 2355 1161 2899 1339
rect 2355 623 2435 1161
rect 2837 953 2899 1161
rect 2729 766 2899 953
rect 2164 558 2435 623
rect 2850 610 2899 766
rect 3029 610 3087 1339
rect 2164 556 2255 558
rect 2850 556 3087 610
rect 421 342 2284 482
rect 421 -158 712 342
rect 1870 -158 2284 342
rect 3337 200 3426 1621
rect 3337 144 3460 200
rect 3337 110 3482 144
rect 4317 110 4377 144
rect 3337 84 4377 110
rect 3337 21 4343 84
rect 421 -185 2284 -158
rect 421 -358 537 -185
rect 421 -374 2284 -358
rect 421 -1094 712 -374
rect 2140 -1094 2284 -374
rect 421 -1188 2284 -1094
rect 2341 -185 4204 -90
rect 2341 -358 2457 -185
rect 2341 -374 4204 -358
rect 2341 -1094 2632 -374
rect 4060 -1094 4204 -374
rect 2341 -1188 4204 -1094
rect 421 -2412 528 -1188
rect 599 -1355 2235 -1266
rect 599 -2470 714 -1355
rect 2120 -2470 2235 -1355
rect 2341 -2028 2448 -1188
rect 2519 -1355 4155 -1266
rect 2519 -2470 2634 -1355
rect 4040 -2470 4155 -1355
rect 471 -2511 4277 -2470
rect 471 -2681 582 -2511
rect 2327 -2681 2502 -2511
rect 4247 -2681 4277 -2511
rect 471 -2743 4277 -2681
rect 387 -2789 421 -2763
rect 4320 -2763 4343 21
rect 4320 -2789 4377 -2763
rect 387 -2823 447 -2789
rect 4317 -2823 4377 -2789
<< viali >>
rect 1221 674 1297 1355
rect 1802 676 1878 1357
rect 2225 623 2355 1352
rect 2899 610 3029 1339
rect 537 -358 2284 -185
rect 2457 -358 4204 -185
rect 582 -2681 2327 -2511
rect 2502 -2681 4247 -2511
<< metal1 >>
rect 393 1541 3150 1563
rect 393 1322 544 1541
rect 842 1357 3150 1541
rect 842 1355 1802 1357
rect 842 1322 1221 1355
rect 393 1306 1221 1322
rect 824 764 888 1306
rect 340 619 540 690
rect 340 567 796 619
rect 888 567 894 619
rect 340 490 540 567
rect 943 411 980 1231
rect 1052 518 1101 1172
rect 1211 674 1221 1306
rect 1297 1306 1802 1355
rect 1297 674 1308 1306
rect 1406 760 1470 1306
rect 1211 659 1308 674
rect 1534 619 1571 1232
rect 1483 567 1489 619
rect 1567 567 1572 619
rect 1052 449 1066 518
rect 1231 449 1245 518
rect 908 330 922 411
rect 1086 330 1099 411
rect 909 200 946 330
rect 1062 200 1099 330
rect 793 138 866 153
rect 793 -46 803 138
rect 857 -46 866 138
rect 793 -59 866 -46
rect 964 -92 1036 156
rect 1158 139 1207 449
rect 1534 401 1571 567
rect 1620 500 1669 1171
rect 1791 676 1802 1306
rect 1878 1352 3150 1357
rect 1878 918 2225 1352
rect 1878 676 1888 918
rect 1791 664 1888 676
rect 2009 619 2080 739
rect 2186 623 2225 918
rect 2355 1339 3150 1352
rect 2355 1201 2899 1339
rect 2355 623 2383 1201
rect 2863 1166 2899 1201
rect 2186 589 2383 623
rect 2009 561 2080 567
rect 1620 451 1792 500
rect 1490 364 1680 401
rect 1490 200 1527 364
rect 1643 200 1680 364
rect 1201 -45 1207 139
rect 1158 -57 1207 -45
rect 1375 140 1448 151
rect 1375 -44 1382 140
rect 1436 -44 1448 140
rect 1375 -61 1448 -44
rect 1552 -92 1624 151
rect 1743 140 1792 451
rect 1786 -44 1792 140
rect 1743 -59 1792 -44
rect 2187 257 2383 589
rect 2446 765 2590 964
rect 2446 221 2497 765
rect 2628 411 2665 1030
rect 2862 954 2899 1166
rect 2729 766 2899 954
rect 2863 610 2899 766
rect 3029 1306 3150 1339
rect 3029 610 3060 1306
rect 2863 577 3060 610
rect 2759 449 2767 518
rect 2951 449 2960 518
rect 2565 330 2576 411
rect 2732 330 2742 411
rect 2879 255 2960 449
rect 2446 150 2592 221
rect 2772 150 2782 221
rect 2879 125 2960 133
rect 2187 -48 2383 -38
rect 2884 -92 2956 -90
rect 3472 -92 3544 -90
rect 326 -185 4398 -92
rect 326 -358 537 -185
rect 2284 -358 2457 -185
rect 4204 -358 4398 -185
rect 326 -368 4398 -358
rect 904 -449 959 -397
rect 1040 -449 1046 -397
rect 904 -453 1046 -449
rect 745 -742 867 -736
rect 745 -895 751 -742
rect 860 -895 867 -742
rect 745 -901 867 -895
rect 904 -1067 939 -453
rect 1370 -455 1376 -402
rect 1457 -455 1525 -402
rect 1370 -458 1525 -455
rect 1190 -501 1292 -495
rect 1190 -685 1196 -501
rect 1286 -685 1292 -501
rect 1190 -691 1292 -685
rect 977 -741 1099 -735
rect 977 -894 984 -741
rect 1093 -894 1099 -741
rect 977 -900 1099 -894
rect 1350 -914 1356 -748
rect 1446 -914 1452 -748
rect 1489 -949 1525 -458
rect 2824 -449 2879 -397
rect 2960 -449 2966 -397
rect 2824 -453 2966 -449
rect 1562 -501 1664 -495
rect 1562 -685 1568 -501
rect 1658 -685 1664 -501
rect 1755 -511 1876 -505
rect 1755 -664 1761 -511
rect 1870 -664 1876 -511
rect 1755 -670 1876 -664
rect 1988 -511 2109 -505
rect 1988 -664 1994 -511
rect 2103 -664 2109 -511
rect 1988 -670 2109 -664
rect 1562 -691 1664 -685
rect 1334 -979 1685 -949
rect 1334 -985 1623 -979
rect 1617 -1039 1623 -985
rect 1679 -1039 1685 -979
rect 1913 -1067 1948 -729
rect 2665 -742 2787 -736
rect 904 -1115 1948 -1067
rect 2209 -953 2393 -776
rect 2665 -895 2671 -742
rect 2780 -895 2787 -742
rect 2665 -901 2787 -895
rect 314 -1168 891 -1164
rect 314 -1368 735 -1168
rect 885 -1368 891 -1168
rect 1051 -1245 1128 -1237
rect 1051 -1307 1128 -1301
rect 1051 -1461 1087 -1307
rect 894 -1489 1087 -1461
rect 1479 -1464 1515 -1115
rect 1728 -1245 1805 -1239
rect 1728 -1309 1805 -1301
rect 887 -1497 1087 -1489
rect 740 -1548 856 -1542
rect 740 -1885 746 -1548
rect 850 -1885 856 -1548
rect 740 -1891 856 -1885
rect 887 -2384 923 -1497
rect 1322 -1500 1515 -1464
rect 1756 -1462 1792 -1309
rect 1756 -1498 1949 -1462
rect 967 -1548 1083 -1542
rect 967 -1885 973 -1548
rect 1077 -1885 1083 -1548
rect 967 -1891 1083 -1885
rect 1323 -1558 1440 -1552
rect 1323 -1882 1329 -1558
rect 1434 -1882 1440 -1558
rect 1323 -1888 1440 -1882
rect 1166 -1987 1282 -1981
rect 1166 -2324 1172 -1987
rect 1276 -2324 1282 -1987
rect 1166 -2330 1282 -2324
rect 1479 -2373 1515 -1500
rect 1552 -1987 1668 -1981
rect 1552 -2324 1558 -1987
rect 1662 -2324 1668 -1987
rect 1552 -2330 1668 -2324
rect 1750 -1987 1866 -1981
rect 1750 -2324 1756 -1987
rect 1860 -2324 1866 -1987
rect 1750 -2330 1866 -2324
rect 1347 -2409 1515 -2373
rect 1910 -2386 1946 -1498
rect 2209 -1826 2217 -953
rect 2387 -1164 2393 -953
rect 2824 -1067 2859 -453
rect 3290 -455 3296 -402
rect 3377 -455 3445 -402
rect 3290 -458 3445 -455
rect 3110 -501 3212 -495
rect 3110 -685 3116 -501
rect 3206 -685 3212 -501
rect 3110 -691 3212 -685
rect 2897 -741 3019 -735
rect 2897 -894 2904 -741
rect 3013 -894 3019 -741
rect 2897 -900 3019 -894
rect 3270 -914 3276 -748
rect 3366 -914 3372 -748
rect 3409 -949 3445 -458
rect 3482 -501 3584 -495
rect 3482 -685 3488 -501
rect 3578 -685 3584 -501
rect 3675 -511 3796 -505
rect 3675 -664 3681 -511
rect 3790 -664 3796 -511
rect 3675 -670 3796 -664
rect 3908 -511 4029 -505
rect 3908 -664 3914 -511
rect 4023 -664 4029 -511
rect 3908 -670 4029 -664
rect 3482 -691 3584 -685
rect 3254 -979 3605 -949
rect 3254 -985 3543 -979
rect 3537 -1039 3543 -985
rect 3599 -1039 3605 -979
rect 3833 -1067 3868 -720
rect 2824 -1115 3868 -1067
rect 4129 -776 4446 -576
rect 4129 -782 4313 -776
rect 2387 -1168 2811 -1164
rect 2387 -1360 2655 -1168
rect 2805 -1360 2811 -1168
rect 2387 -1364 2811 -1360
rect 2971 -1245 3048 -1237
rect 2971 -1307 3048 -1301
rect 2387 -1826 2393 -1364
rect 2971 -1461 3007 -1307
rect 2814 -1489 3007 -1461
rect 3399 -1464 3435 -1115
rect 3648 -1245 3725 -1239
rect 3648 -1309 3725 -1301
rect 2807 -1497 3007 -1489
rect 2209 -1836 2393 -1826
rect 2660 -1548 2776 -1542
rect 2660 -1885 2666 -1548
rect 2770 -1885 2776 -1548
rect 2660 -1891 2776 -1885
rect 1978 -1987 2094 -1981
rect 1978 -2324 1984 -1987
rect 2088 -2324 2094 -1987
rect 1978 -2330 2094 -2324
rect 2807 -2384 2843 -1497
rect 3242 -1500 3435 -1464
rect 3676 -1462 3712 -1309
rect 3676 -1498 3869 -1462
rect 2887 -1548 3003 -1542
rect 2887 -1885 2893 -1548
rect 2997 -1885 3003 -1548
rect 2887 -1891 3003 -1885
rect 3243 -1558 3360 -1552
rect 3243 -1882 3249 -1558
rect 3354 -1882 3360 -1558
rect 3243 -1888 3360 -1882
rect 3086 -1987 3202 -1981
rect 3086 -2324 3092 -1987
rect 3196 -2324 3202 -1987
rect 3086 -2330 3202 -2324
rect 3399 -2373 3435 -1500
rect 3472 -1987 3588 -1981
rect 3472 -2324 3478 -1987
rect 3582 -2324 3588 -1987
rect 3472 -2330 3588 -2324
rect 3670 -1987 3786 -1981
rect 3670 -2324 3676 -1987
rect 3780 -2324 3786 -1987
rect 3670 -2330 3786 -2324
rect 3267 -2409 3435 -2373
rect 3830 -2386 3866 -1498
rect 4129 -1826 4137 -782
rect 4307 -1826 4313 -782
rect 4129 -1836 4313 -1826
rect 3898 -1987 4014 -1981
rect 3898 -2324 3904 -1987
rect 4008 -2324 4014 -1987
rect 3898 -2330 4014 -2324
rect 328 -2479 4435 -2470
rect 328 -2698 542 -2479
rect 840 -2511 2462 -2479
rect 2760 -2511 4435 -2479
rect 2327 -2681 2462 -2511
rect 4247 -2681 4435 -2511
rect 840 -2698 2462 -2681
rect 2760 -2698 4435 -2681
rect 328 -2705 4435 -2698
<< via1 >>
rect 544 1322 842 1541
rect 796 567 888 619
rect 1489 567 1567 619
rect 1066 449 1231 518
rect 922 330 1086 411
rect 803 -46 857 138
rect 2009 567 2080 619
rect 1147 -45 1201 139
rect 1382 -44 1436 140
rect 1732 -44 1786 140
rect 2187 -38 2383 257
rect 2767 449 2951 518
rect 2576 330 2732 411
rect 2592 150 2772 221
rect 2879 133 2960 255
rect 959 -449 1040 -397
rect 751 -895 860 -742
rect 1376 -455 1457 -402
rect 1196 -685 1286 -501
rect 984 -894 1093 -741
rect 1356 -914 1446 -748
rect 2879 -449 2960 -397
rect 1568 -685 1658 -501
rect 1761 -664 1870 -511
rect 1994 -664 2103 -511
rect 1623 -1039 1679 -979
rect 2671 -895 2780 -742
rect 735 -1368 885 -1168
rect 1051 -1301 1128 -1245
rect 1728 -1301 1805 -1245
rect 746 -1885 850 -1548
rect 973 -1885 1077 -1548
rect 1329 -1882 1434 -1558
rect 1172 -2324 1276 -1987
rect 1558 -2324 1662 -1987
rect 1756 -2324 1860 -1987
rect 2217 -1826 2387 -953
rect 3296 -455 3377 -402
rect 3116 -685 3206 -501
rect 2904 -894 3013 -741
rect 3276 -914 3366 -748
rect 3488 -685 3578 -501
rect 3681 -664 3790 -511
rect 3914 -664 4023 -511
rect 3543 -1039 3599 -979
rect 2655 -1360 2805 -1168
rect 2971 -1301 3048 -1245
rect 3648 -1301 3725 -1245
rect 2666 -1885 2770 -1548
rect 1984 -2324 2088 -1987
rect 2893 -1885 2997 -1548
rect 3249 -1882 3354 -1558
rect 3092 -2324 3196 -1987
rect 3478 -2324 3582 -1987
rect 3676 -2324 3780 -1987
rect 4137 -1826 4307 -782
rect 3904 -2324 4008 -1987
rect 542 -2511 840 -2479
rect 2462 -2511 2760 -2479
rect 542 -2681 582 -2511
rect 582 -2681 840 -2511
rect 2462 -2681 2502 -2511
rect 2502 -2681 2760 -2511
rect 542 -2698 840 -2681
rect 2462 -2698 2760 -2681
<< metal2 >>
rect 529 1541 867 1556
rect 529 1322 544 1541
rect 842 1322 867 1541
rect 529 1306 867 1322
rect 529 -2470 660 1306
rect 789 567 796 619
rect 888 567 1489 619
rect 1567 567 2009 619
rect 2080 567 2087 619
rect 1052 449 1066 518
rect 1231 449 2767 518
rect 2951 449 2960 518
rect 908 330 922 411
rect 1086 330 2576 411
rect 2732 330 3377 411
rect 1376 142 1457 330
rect 2187 257 2383 269
rect 795 139 1207 141
rect 795 138 1147 139
rect 795 -46 803 138
rect 857 -45 1147 138
rect 1201 -45 1207 139
rect 857 -46 1207 -45
rect 795 -47 1207 -46
rect 1376 140 1792 142
rect 1376 -44 1382 140
rect 1436 -44 1732 140
rect 1786 -44 1792 140
rect 1376 -46 1792 -44
rect 2879 255 2960 263
rect 2579 150 2592 221
rect 2772 150 2782 221
rect 959 -397 1040 -47
rect 959 -455 1040 -449
rect 1376 -402 1457 -46
rect 2187 -90 2383 -38
rect 2187 -382 2580 -90
rect 1376 -461 1457 -455
rect 736 -501 2393 -489
rect 736 -685 1196 -501
rect 1286 -685 1568 -501
rect 1658 -511 2393 -501
rect 1658 -664 1761 -511
rect 1870 -664 1994 -511
rect 2103 -664 2393 -511
rect 1658 -685 2393 -664
rect 736 -693 2393 -685
rect 732 -741 2127 -734
rect 732 -742 984 -741
rect 732 -895 751 -742
rect 860 -894 984 -742
rect 1093 -748 2127 -741
rect 1093 -894 1356 -748
rect 860 -895 1356 -894
rect 732 -914 1356 -895
rect 1446 -914 2127 -748
rect 732 -938 2127 -914
rect 732 -1168 891 -938
rect 2209 -953 2393 -693
rect 732 -1368 735 -1168
rect 885 -1368 891 -1168
rect 1623 -979 1679 -972
rect 1623 -1245 1679 -1039
rect 1043 -1301 1051 -1245
rect 1128 -1301 1728 -1245
rect 1805 -1301 1816 -1245
rect 732 -1513 891 -1368
rect 732 -1548 2122 -1513
rect 732 -1885 746 -1548
rect 850 -1885 973 -1548
rect 1077 -1558 2122 -1548
rect 1077 -1882 1329 -1558
rect 1434 -1882 2122 -1558
rect 1077 -1885 2122 -1882
rect 732 -1897 2122 -1885
rect 2209 -1826 2217 -953
rect 2387 -1826 2393 -953
rect 2209 -1958 2393 -1826
rect 733 -1987 2393 -1958
rect 733 -2324 1172 -1987
rect 1276 -2324 1558 -1987
rect 1662 -2324 1756 -1987
rect 1860 -2324 1984 -1987
rect 2088 -2324 2393 -1987
rect 733 -2342 2393 -2324
rect 2449 -2470 2580 -382
rect 2653 -734 2715 150
rect 2879 -397 2960 133
rect 2879 -455 2960 -449
rect 3296 -402 3377 330
rect 3296 -461 3377 -455
rect 2761 -501 4313 -489
rect 2761 -685 3116 -501
rect 3206 -685 3488 -501
rect 3578 -511 4313 -501
rect 3578 -664 3681 -511
rect 3790 -664 3914 -511
rect 4023 -664 4313 -511
rect 3578 -685 4313 -664
rect 2761 -693 4313 -685
rect 2652 -741 4047 -734
rect 2652 -742 2904 -741
rect 2652 -895 2671 -742
rect 2780 -894 2904 -742
rect 3013 -748 4047 -741
rect 3013 -894 3276 -748
rect 2780 -895 3276 -894
rect 2652 -914 3276 -895
rect 3366 -914 4047 -748
rect 2652 -938 4047 -914
rect 4129 -782 4313 -693
rect 2652 -1168 2811 -938
rect 2652 -1360 2655 -1168
rect 2805 -1360 2811 -1168
rect 3543 -979 3599 -972
rect 3543 -1245 3599 -1039
rect 2963 -1301 2971 -1245
rect 3048 -1301 3648 -1245
rect 3725 -1301 3736 -1245
rect 2652 -1513 2811 -1360
rect 2652 -1548 4042 -1513
rect 2652 -1885 2666 -1548
rect 2770 -1885 2893 -1548
rect 2997 -1558 4042 -1548
rect 2997 -1882 3249 -1558
rect 3354 -1882 4042 -1558
rect 2997 -1885 4042 -1882
rect 2652 -1897 4042 -1885
rect 4129 -1826 4137 -782
rect 4307 -1826 4313 -782
rect 4129 -1958 4313 -1826
rect 2653 -1987 4313 -1958
rect 2653 -2324 3092 -1987
rect 3196 -2324 3478 -1987
rect 3582 -2324 3676 -1987
rect 3780 -2324 3904 -1987
rect 4008 -2324 4313 -1987
rect 2653 -2342 4313 -2324
rect 529 -2479 849 -2470
rect 529 -2698 542 -2479
rect 840 -2698 849 -2479
rect 529 -2705 849 -2698
rect 2449 -2479 2769 -2470
rect 2449 -2698 2462 -2479
rect 2760 -2698 2769 -2479
rect 2449 -2705 2769 -2698
use sky130_fd_pr__nfet_g5v0d10v5_HRGQF2  sky130_fd_pr__nfet_g5v0d10v5_HRGQF2_0 paramcells
timestamp 1713821214
transform -1 0 3337 0 1 -1936
box -357 -658 357 658
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4  sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4_0 paramcells
timestamp 1713821214
transform -1 0 2828 0 1 -1935
box -278 -658 278 658
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4  sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4_1
timestamp 1713821214
transform 1 0 3848 0 1 -1935
box -278 -658 278 658
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ3N  sky130_fd_pr__nfet_g5v0d10v5_UNEQ3N_0 paramcells
timestamp 1713820565
transform 1 0 2647 0 -1 867
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6  sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6_0 paramcells
timestamp 1713821214
transform 1 0 3347 0 1 -738
box -387 -462 387 462
use sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6  sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_0 paramcells
timestamp 1713821214
transform 1 0 922 0 1 -738
box -308 -462 308 462
use sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6  sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_1
timestamp 1713821214
transform 1 0 2842 0 1 -738
box -308 -462 308 462
use sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6  sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_2
timestamp 1713821214
transform 1 0 3852 0 1 -738
box -308 -462 308 462
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 paramcells
timestamp 1652924542
transform 1 0 1585 0 -1 82
box -387 -362 387 362
use sky130_fd_pr__diode_pw2nd_05v5_FT76RK  XD1 paramcells
timestamp 1713888873
transform 1 0 2045 0 -1 703
box -183 -183 183 183
use sky130_fd_pr__nfet_g5v0d10v5_HRGQF2  XM1
timestamp 1713821214
transform -1 0 1417 0 1 -1936
box -357 -658 357 658
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4  XM3
timestamp 1713821214
transform -1 0 908 0 1 -1935
box -278 -658 278 658
use sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6  XM4
timestamp 1713821214
transform 1 0 1427 0 1 -738
box -387 -462 387 462
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4  XM5
timestamp 1713821214
transform 1 0 1928 0 1 -1935
box -278 -658 278 658
use sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6  XM6
timestamp 1713821214
transform 1 0 1932 0 1 -738
box -308 -462 308 462
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM7
timestamp 1652924542
transform 1 0 1001 0 -1 82
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM8 paramcells
timestamp 1652200182
transform 1 0 964 0 -1 966
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM10
timestamp 1652200182
transform 1 0 1546 0 -1 966
box -278 -458 278 458
<< labels >>
flabel metal1 326 -352 526 -152 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 4246 -776 4446 -576 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 340 490 540 690 0 FreeSans 256 0 0 0 on
port 1 nsew
flabel metal1 1705 473 1705 473 0 FreeSans 320 0 0 0 onb
flabel metal1 1068 647 1068 647 0 FreeSans 320 0 0 0 onp
flabel metal1 314 -1364 514 -1164 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 336 -2691 536 -2491 0 FreeSans 256 0 0 0 vss
port 2 nsew
<< end >>
