magic
tech sky130A
magscale 1 2
timestamp 1713888873
<< pwell >>
rect -2779 -558 2779 558
<< mvnnmos >>
rect -2551 -300 -2351 300
rect -2293 -300 -2093 300
rect -2035 -300 -1835 300
rect -1777 -300 -1577 300
rect -1519 -300 -1319 300
rect -1261 -300 -1061 300
rect -1003 -300 -803 300
rect -745 -300 -545 300
rect -487 -300 -287 300
rect -229 -300 -29 300
rect 29 -300 229 300
rect 287 -300 487 300
rect 545 -300 745 300
rect 803 -300 1003 300
rect 1061 -300 1261 300
rect 1319 -300 1519 300
rect 1577 -300 1777 300
rect 1835 -300 2035 300
rect 2093 -300 2293 300
rect 2351 -300 2551 300
<< mvndiff >>
rect -2609 288 -2551 300
rect -2609 -288 -2597 288
rect -2563 -288 -2551 288
rect -2609 -300 -2551 -288
rect -2351 288 -2293 300
rect -2351 -288 -2339 288
rect -2305 -288 -2293 288
rect -2351 -300 -2293 -288
rect -2093 288 -2035 300
rect -2093 -288 -2081 288
rect -2047 -288 -2035 288
rect -2093 -300 -2035 -288
rect -1835 288 -1777 300
rect -1835 -288 -1823 288
rect -1789 -288 -1777 288
rect -1835 -300 -1777 -288
rect -1577 288 -1519 300
rect -1577 -288 -1565 288
rect -1531 -288 -1519 288
rect -1577 -300 -1519 -288
rect -1319 288 -1261 300
rect -1319 -288 -1307 288
rect -1273 -288 -1261 288
rect -1319 -300 -1261 -288
rect -1061 288 -1003 300
rect -1061 -288 -1049 288
rect -1015 -288 -1003 288
rect -1061 -300 -1003 -288
rect -803 288 -745 300
rect -803 -288 -791 288
rect -757 -288 -745 288
rect -803 -300 -745 -288
rect -545 288 -487 300
rect -545 -288 -533 288
rect -499 -288 -487 288
rect -545 -300 -487 -288
rect -287 288 -229 300
rect -287 -288 -275 288
rect -241 -288 -229 288
rect -287 -300 -229 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 229 288 287 300
rect 229 -288 241 288
rect 275 -288 287 288
rect 229 -300 287 -288
rect 487 288 545 300
rect 487 -288 499 288
rect 533 -288 545 288
rect 487 -300 545 -288
rect 745 288 803 300
rect 745 -288 757 288
rect 791 -288 803 288
rect 745 -300 803 -288
rect 1003 288 1061 300
rect 1003 -288 1015 288
rect 1049 -288 1061 288
rect 1003 -300 1061 -288
rect 1261 288 1319 300
rect 1261 -288 1273 288
rect 1307 -288 1319 288
rect 1261 -300 1319 -288
rect 1519 288 1577 300
rect 1519 -288 1531 288
rect 1565 -288 1577 288
rect 1519 -300 1577 -288
rect 1777 288 1835 300
rect 1777 -288 1789 288
rect 1823 -288 1835 288
rect 1777 -300 1835 -288
rect 2035 288 2093 300
rect 2035 -288 2047 288
rect 2081 -288 2093 288
rect 2035 -300 2093 -288
rect 2293 288 2351 300
rect 2293 -288 2305 288
rect 2339 -288 2351 288
rect 2293 -300 2351 -288
rect 2551 288 2609 300
rect 2551 -288 2563 288
rect 2597 -288 2609 288
rect 2551 -300 2609 -288
<< mvndiffc >>
rect -2597 -288 -2563 288
rect -2339 -288 -2305 288
rect -2081 -288 -2047 288
rect -1823 -288 -1789 288
rect -1565 -288 -1531 288
rect -1307 -288 -1273 288
rect -1049 -288 -1015 288
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect 1015 -288 1049 288
rect 1273 -288 1307 288
rect 1531 -288 1565 288
rect 1789 -288 1823 288
rect 2047 -288 2081 288
rect 2305 -288 2339 288
rect 2563 -288 2597 288
<< mvpsubdiff >>
rect -2743 510 2743 522
rect -2743 476 -2635 510
rect 2635 476 2743 510
rect -2743 464 2743 476
rect -2743 414 -2685 464
rect -2743 -414 -2731 414
rect -2697 -414 -2685 414
rect 2685 414 2743 464
rect -2743 -464 -2685 -414
rect 2685 -414 2697 414
rect 2731 -414 2743 414
rect 2685 -464 2743 -414
rect -2743 -476 2743 -464
rect -2743 -510 -2635 -476
rect 2635 -510 2743 -476
rect -2743 -522 2743 -510
<< mvpsubdiffcont >>
rect -2635 476 2635 510
rect -2731 -414 -2697 414
rect 2697 -414 2731 414
rect -2635 -510 2635 -476
<< poly >>
rect -2551 372 -2351 388
rect -2551 338 -2535 372
rect -2367 338 -2351 372
rect -2551 300 -2351 338
rect -2293 372 -2093 388
rect -2293 338 -2277 372
rect -2109 338 -2093 372
rect -2293 300 -2093 338
rect -2035 372 -1835 388
rect -2035 338 -2019 372
rect -1851 338 -1835 372
rect -2035 300 -1835 338
rect -1777 372 -1577 388
rect -1777 338 -1761 372
rect -1593 338 -1577 372
rect -1777 300 -1577 338
rect -1519 372 -1319 388
rect -1519 338 -1503 372
rect -1335 338 -1319 372
rect -1519 300 -1319 338
rect -1261 372 -1061 388
rect -1261 338 -1245 372
rect -1077 338 -1061 372
rect -1261 300 -1061 338
rect -1003 372 -803 388
rect -1003 338 -987 372
rect -819 338 -803 372
rect -1003 300 -803 338
rect -745 372 -545 388
rect -745 338 -729 372
rect -561 338 -545 372
rect -745 300 -545 338
rect -487 372 -287 388
rect -487 338 -471 372
rect -303 338 -287 372
rect -487 300 -287 338
rect -229 372 -29 388
rect -229 338 -213 372
rect -45 338 -29 372
rect -229 300 -29 338
rect 29 372 229 388
rect 29 338 45 372
rect 213 338 229 372
rect 29 300 229 338
rect 287 372 487 388
rect 287 338 303 372
rect 471 338 487 372
rect 287 300 487 338
rect 545 372 745 388
rect 545 338 561 372
rect 729 338 745 372
rect 545 300 745 338
rect 803 372 1003 388
rect 803 338 819 372
rect 987 338 1003 372
rect 803 300 1003 338
rect 1061 372 1261 388
rect 1061 338 1077 372
rect 1245 338 1261 372
rect 1061 300 1261 338
rect 1319 372 1519 388
rect 1319 338 1335 372
rect 1503 338 1519 372
rect 1319 300 1519 338
rect 1577 372 1777 388
rect 1577 338 1593 372
rect 1761 338 1777 372
rect 1577 300 1777 338
rect 1835 372 2035 388
rect 1835 338 1851 372
rect 2019 338 2035 372
rect 1835 300 2035 338
rect 2093 372 2293 388
rect 2093 338 2109 372
rect 2277 338 2293 372
rect 2093 300 2293 338
rect 2351 372 2551 388
rect 2351 338 2367 372
rect 2535 338 2551 372
rect 2351 300 2551 338
rect -2551 -338 -2351 -300
rect -2551 -372 -2535 -338
rect -2367 -372 -2351 -338
rect -2551 -388 -2351 -372
rect -2293 -338 -2093 -300
rect -2293 -372 -2277 -338
rect -2109 -372 -2093 -338
rect -2293 -388 -2093 -372
rect -2035 -338 -1835 -300
rect -2035 -372 -2019 -338
rect -1851 -372 -1835 -338
rect -2035 -388 -1835 -372
rect -1777 -338 -1577 -300
rect -1777 -372 -1761 -338
rect -1593 -372 -1577 -338
rect -1777 -388 -1577 -372
rect -1519 -338 -1319 -300
rect -1519 -372 -1503 -338
rect -1335 -372 -1319 -338
rect -1519 -388 -1319 -372
rect -1261 -338 -1061 -300
rect -1261 -372 -1245 -338
rect -1077 -372 -1061 -338
rect -1261 -388 -1061 -372
rect -1003 -338 -803 -300
rect -1003 -372 -987 -338
rect -819 -372 -803 -338
rect -1003 -388 -803 -372
rect -745 -338 -545 -300
rect -745 -372 -729 -338
rect -561 -372 -545 -338
rect -745 -388 -545 -372
rect -487 -338 -287 -300
rect -487 -372 -471 -338
rect -303 -372 -287 -338
rect -487 -388 -287 -372
rect -229 -338 -29 -300
rect -229 -372 -213 -338
rect -45 -372 -29 -338
rect -229 -388 -29 -372
rect 29 -338 229 -300
rect 29 -372 45 -338
rect 213 -372 229 -338
rect 29 -388 229 -372
rect 287 -338 487 -300
rect 287 -372 303 -338
rect 471 -372 487 -338
rect 287 -388 487 -372
rect 545 -338 745 -300
rect 545 -372 561 -338
rect 729 -372 745 -338
rect 545 -388 745 -372
rect 803 -338 1003 -300
rect 803 -372 819 -338
rect 987 -372 1003 -338
rect 803 -388 1003 -372
rect 1061 -338 1261 -300
rect 1061 -372 1077 -338
rect 1245 -372 1261 -338
rect 1061 -388 1261 -372
rect 1319 -338 1519 -300
rect 1319 -372 1335 -338
rect 1503 -372 1519 -338
rect 1319 -388 1519 -372
rect 1577 -338 1777 -300
rect 1577 -372 1593 -338
rect 1761 -372 1777 -338
rect 1577 -388 1777 -372
rect 1835 -338 2035 -300
rect 1835 -372 1851 -338
rect 2019 -372 2035 -338
rect 1835 -388 2035 -372
rect 2093 -338 2293 -300
rect 2093 -372 2109 -338
rect 2277 -372 2293 -338
rect 2093 -388 2293 -372
rect 2351 -338 2551 -300
rect 2351 -372 2367 -338
rect 2535 -372 2551 -338
rect 2351 -388 2551 -372
<< polycont >>
rect -2535 338 -2367 372
rect -2277 338 -2109 372
rect -2019 338 -1851 372
rect -1761 338 -1593 372
rect -1503 338 -1335 372
rect -1245 338 -1077 372
rect -987 338 -819 372
rect -729 338 -561 372
rect -471 338 -303 372
rect -213 338 -45 372
rect 45 338 213 372
rect 303 338 471 372
rect 561 338 729 372
rect 819 338 987 372
rect 1077 338 1245 372
rect 1335 338 1503 372
rect 1593 338 1761 372
rect 1851 338 2019 372
rect 2109 338 2277 372
rect 2367 338 2535 372
rect -2535 -372 -2367 -338
rect -2277 -372 -2109 -338
rect -2019 -372 -1851 -338
rect -1761 -372 -1593 -338
rect -1503 -372 -1335 -338
rect -1245 -372 -1077 -338
rect -987 -372 -819 -338
rect -729 -372 -561 -338
rect -471 -372 -303 -338
rect -213 -372 -45 -338
rect 45 -372 213 -338
rect 303 -372 471 -338
rect 561 -372 729 -338
rect 819 -372 987 -338
rect 1077 -372 1245 -338
rect 1335 -372 1503 -338
rect 1593 -372 1761 -338
rect 1851 -372 2019 -338
rect 2109 -372 2277 -338
rect 2367 -372 2535 -338
<< locali >>
rect -2731 476 -2635 510
rect 2635 476 2731 510
rect -2731 414 -2697 476
rect 2697 414 2731 476
rect -2551 338 -2535 372
rect -2367 338 -2351 372
rect -2293 338 -2277 372
rect -2109 338 -2093 372
rect -2035 338 -2019 372
rect -1851 338 -1835 372
rect -1777 338 -1761 372
rect -1593 338 -1577 372
rect -1519 338 -1503 372
rect -1335 338 -1319 372
rect -1261 338 -1245 372
rect -1077 338 -1061 372
rect -1003 338 -987 372
rect -819 338 -803 372
rect -745 338 -729 372
rect -561 338 -545 372
rect -487 338 -471 372
rect -303 338 -287 372
rect -229 338 -213 372
rect -45 338 -29 372
rect 29 338 45 372
rect 213 338 229 372
rect 287 338 303 372
rect 471 338 487 372
rect 545 338 561 372
rect 729 338 745 372
rect 803 338 819 372
rect 987 338 1003 372
rect 1061 338 1077 372
rect 1245 338 1261 372
rect 1319 338 1335 372
rect 1503 338 1519 372
rect 1577 338 1593 372
rect 1761 338 1777 372
rect 1835 338 1851 372
rect 2019 338 2035 372
rect 2093 338 2109 372
rect 2277 338 2293 372
rect 2351 338 2367 372
rect 2535 338 2551 372
rect -2597 288 -2563 304
rect -2597 -304 -2563 -288
rect -2339 288 -2305 304
rect -2339 -304 -2305 -288
rect -2081 288 -2047 304
rect -2081 -304 -2047 -288
rect -1823 288 -1789 304
rect -1823 -304 -1789 -288
rect -1565 288 -1531 304
rect -1565 -304 -1531 -288
rect -1307 288 -1273 304
rect -1307 -304 -1273 -288
rect -1049 288 -1015 304
rect -1049 -304 -1015 -288
rect -791 288 -757 304
rect -791 -304 -757 -288
rect -533 288 -499 304
rect -533 -304 -499 -288
rect -275 288 -241 304
rect -275 -304 -241 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 241 288 275 304
rect 241 -304 275 -288
rect 499 288 533 304
rect 499 -304 533 -288
rect 757 288 791 304
rect 757 -304 791 -288
rect 1015 288 1049 304
rect 1015 -304 1049 -288
rect 1273 288 1307 304
rect 1273 -304 1307 -288
rect 1531 288 1565 304
rect 1531 -304 1565 -288
rect 1789 288 1823 304
rect 1789 -304 1823 -288
rect 2047 288 2081 304
rect 2047 -304 2081 -288
rect 2305 288 2339 304
rect 2305 -304 2339 -288
rect 2563 288 2597 304
rect 2563 -304 2597 -288
rect -2551 -372 -2535 -338
rect -2367 -372 -2351 -338
rect -2293 -372 -2277 -338
rect -2109 -372 -2093 -338
rect -2035 -372 -2019 -338
rect -1851 -372 -1835 -338
rect -1777 -372 -1761 -338
rect -1593 -372 -1577 -338
rect -1519 -372 -1503 -338
rect -1335 -372 -1319 -338
rect -1261 -372 -1245 -338
rect -1077 -372 -1061 -338
rect -1003 -372 -987 -338
rect -819 -372 -803 -338
rect -745 -372 -729 -338
rect -561 -372 -545 -338
rect -487 -372 -471 -338
rect -303 -372 -287 -338
rect -229 -372 -213 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 213 -372 229 -338
rect 287 -372 303 -338
rect 471 -372 487 -338
rect 545 -372 561 -338
rect 729 -372 745 -338
rect 803 -372 819 -338
rect 987 -372 1003 -338
rect 1061 -372 1077 -338
rect 1245 -372 1261 -338
rect 1319 -372 1335 -338
rect 1503 -372 1519 -338
rect 1577 -372 1593 -338
rect 1761 -372 1777 -338
rect 1835 -372 1851 -338
rect 2019 -372 2035 -338
rect 2093 -372 2109 -338
rect 2277 -372 2293 -338
rect 2351 -372 2367 -338
rect 2535 -372 2551 -338
rect -2731 -476 -2697 -414
rect 2697 -476 2731 -414
rect -2731 -510 -2635 -476
rect 2635 -510 2731 -476
<< viali >>
rect -2535 338 -2367 372
rect -2277 338 -2109 372
rect -2019 338 -1851 372
rect -1761 338 -1593 372
rect -1503 338 -1335 372
rect -1245 338 -1077 372
rect -987 338 -819 372
rect -729 338 -561 372
rect -471 338 -303 372
rect -213 338 -45 372
rect 45 338 213 372
rect 303 338 471 372
rect 561 338 729 372
rect 819 338 987 372
rect 1077 338 1245 372
rect 1335 338 1503 372
rect 1593 338 1761 372
rect 1851 338 2019 372
rect 2109 338 2277 372
rect 2367 338 2535 372
rect -2597 -288 -2563 288
rect -2339 -288 -2305 288
rect -2081 -288 -2047 288
rect -1823 -288 -1789 288
rect -1565 -288 -1531 288
rect -1307 -288 -1273 288
rect -1049 -288 -1015 288
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect 1015 -288 1049 288
rect 1273 -288 1307 288
rect 1531 -288 1565 288
rect 1789 -288 1823 288
rect 2047 -288 2081 288
rect 2305 -288 2339 288
rect 2563 -288 2597 288
rect -2535 -372 -2367 -338
rect -2277 -372 -2109 -338
rect -2019 -372 -1851 -338
rect -1761 -372 -1593 -338
rect -1503 -372 -1335 -338
rect -1245 -372 -1077 -338
rect -987 -372 -819 -338
rect -729 -372 -561 -338
rect -471 -372 -303 -338
rect -213 -372 -45 -338
rect 45 -372 213 -338
rect 303 -372 471 -338
rect 561 -372 729 -338
rect 819 -372 987 -338
rect 1077 -372 1245 -338
rect 1335 -372 1503 -338
rect 1593 -372 1761 -338
rect 1851 -372 2019 -338
rect 2109 -372 2277 -338
rect 2367 -372 2535 -338
<< metal1 >>
rect -2547 372 -2355 378
rect -2547 338 -2535 372
rect -2367 338 -2355 372
rect -2547 332 -2355 338
rect -2289 372 -2097 378
rect -2289 338 -2277 372
rect -2109 338 -2097 372
rect -2289 332 -2097 338
rect -2031 372 -1839 378
rect -2031 338 -2019 372
rect -1851 338 -1839 372
rect -2031 332 -1839 338
rect -1773 372 -1581 378
rect -1773 338 -1761 372
rect -1593 338 -1581 372
rect -1773 332 -1581 338
rect -1515 372 -1323 378
rect -1515 338 -1503 372
rect -1335 338 -1323 372
rect -1515 332 -1323 338
rect -1257 372 -1065 378
rect -1257 338 -1245 372
rect -1077 338 -1065 372
rect -1257 332 -1065 338
rect -999 372 -807 378
rect -999 338 -987 372
rect -819 338 -807 372
rect -999 332 -807 338
rect -741 372 -549 378
rect -741 338 -729 372
rect -561 338 -549 372
rect -741 332 -549 338
rect -483 372 -291 378
rect -483 338 -471 372
rect -303 338 -291 372
rect -483 332 -291 338
rect -225 372 -33 378
rect -225 338 -213 372
rect -45 338 -33 372
rect -225 332 -33 338
rect 33 372 225 378
rect 33 338 45 372
rect 213 338 225 372
rect 33 332 225 338
rect 291 372 483 378
rect 291 338 303 372
rect 471 338 483 372
rect 291 332 483 338
rect 549 372 741 378
rect 549 338 561 372
rect 729 338 741 372
rect 549 332 741 338
rect 807 372 999 378
rect 807 338 819 372
rect 987 338 999 372
rect 807 332 999 338
rect 1065 372 1257 378
rect 1065 338 1077 372
rect 1245 338 1257 372
rect 1065 332 1257 338
rect 1323 372 1515 378
rect 1323 338 1335 372
rect 1503 338 1515 372
rect 1323 332 1515 338
rect 1581 372 1773 378
rect 1581 338 1593 372
rect 1761 338 1773 372
rect 1581 332 1773 338
rect 1839 372 2031 378
rect 1839 338 1851 372
rect 2019 338 2031 372
rect 1839 332 2031 338
rect 2097 372 2289 378
rect 2097 338 2109 372
rect 2277 338 2289 372
rect 2097 332 2289 338
rect 2355 372 2547 378
rect 2355 338 2367 372
rect 2535 338 2547 372
rect 2355 332 2547 338
rect -2603 288 -2557 300
rect -2603 -288 -2597 288
rect -2563 -288 -2557 288
rect -2603 -300 -2557 -288
rect -2345 288 -2299 300
rect -2345 -288 -2339 288
rect -2305 -288 -2299 288
rect -2345 -300 -2299 -288
rect -2087 288 -2041 300
rect -2087 -288 -2081 288
rect -2047 -288 -2041 288
rect -2087 -300 -2041 -288
rect -1829 288 -1783 300
rect -1829 -288 -1823 288
rect -1789 -288 -1783 288
rect -1829 -300 -1783 -288
rect -1571 288 -1525 300
rect -1571 -288 -1565 288
rect -1531 -288 -1525 288
rect -1571 -300 -1525 -288
rect -1313 288 -1267 300
rect -1313 -288 -1307 288
rect -1273 -288 -1267 288
rect -1313 -300 -1267 -288
rect -1055 288 -1009 300
rect -1055 -288 -1049 288
rect -1015 -288 -1009 288
rect -1055 -300 -1009 -288
rect -797 288 -751 300
rect -797 -288 -791 288
rect -757 -288 -751 288
rect -797 -300 -751 -288
rect -539 288 -493 300
rect -539 -288 -533 288
rect -499 -288 -493 288
rect -539 -300 -493 -288
rect -281 288 -235 300
rect -281 -288 -275 288
rect -241 -288 -235 288
rect -281 -300 -235 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 235 288 281 300
rect 235 -288 241 288
rect 275 -288 281 288
rect 235 -300 281 -288
rect 493 288 539 300
rect 493 -288 499 288
rect 533 -288 539 288
rect 493 -300 539 -288
rect 751 288 797 300
rect 751 -288 757 288
rect 791 -288 797 288
rect 751 -300 797 -288
rect 1009 288 1055 300
rect 1009 -288 1015 288
rect 1049 -288 1055 288
rect 1009 -300 1055 -288
rect 1267 288 1313 300
rect 1267 -288 1273 288
rect 1307 -288 1313 288
rect 1267 -300 1313 -288
rect 1525 288 1571 300
rect 1525 -288 1531 288
rect 1565 -288 1571 288
rect 1525 -300 1571 -288
rect 1783 288 1829 300
rect 1783 -288 1789 288
rect 1823 -288 1829 288
rect 1783 -300 1829 -288
rect 2041 288 2087 300
rect 2041 -288 2047 288
rect 2081 -288 2087 288
rect 2041 -300 2087 -288
rect 2299 288 2345 300
rect 2299 -288 2305 288
rect 2339 -288 2345 288
rect 2299 -300 2345 -288
rect 2557 288 2603 300
rect 2557 -288 2563 288
rect 2597 -288 2603 288
rect 2557 -300 2603 -288
rect -2547 -338 -2355 -332
rect -2547 -372 -2535 -338
rect -2367 -372 -2355 -338
rect -2547 -378 -2355 -372
rect -2289 -338 -2097 -332
rect -2289 -372 -2277 -338
rect -2109 -372 -2097 -338
rect -2289 -378 -2097 -372
rect -2031 -338 -1839 -332
rect -2031 -372 -2019 -338
rect -1851 -372 -1839 -338
rect -2031 -378 -1839 -372
rect -1773 -338 -1581 -332
rect -1773 -372 -1761 -338
rect -1593 -372 -1581 -338
rect -1773 -378 -1581 -372
rect -1515 -338 -1323 -332
rect -1515 -372 -1503 -338
rect -1335 -372 -1323 -338
rect -1515 -378 -1323 -372
rect -1257 -338 -1065 -332
rect -1257 -372 -1245 -338
rect -1077 -372 -1065 -338
rect -1257 -378 -1065 -372
rect -999 -338 -807 -332
rect -999 -372 -987 -338
rect -819 -372 -807 -338
rect -999 -378 -807 -372
rect -741 -338 -549 -332
rect -741 -372 -729 -338
rect -561 -372 -549 -338
rect -741 -378 -549 -372
rect -483 -338 -291 -332
rect -483 -372 -471 -338
rect -303 -372 -291 -338
rect -483 -378 -291 -372
rect -225 -338 -33 -332
rect -225 -372 -213 -338
rect -45 -372 -33 -338
rect -225 -378 -33 -372
rect 33 -338 225 -332
rect 33 -372 45 -338
rect 213 -372 225 -338
rect 33 -378 225 -372
rect 291 -338 483 -332
rect 291 -372 303 -338
rect 471 -372 483 -338
rect 291 -378 483 -372
rect 549 -338 741 -332
rect 549 -372 561 -338
rect 729 -372 741 -338
rect 549 -378 741 -372
rect 807 -338 999 -332
rect 807 -372 819 -338
rect 987 -372 999 -338
rect 807 -378 999 -372
rect 1065 -338 1257 -332
rect 1065 -372 1077 -338
rect 1245 -372 1257 -338
rect 1065 -378 1257 -372
rect 1323 -338 1515 -332
rect 1323 -372 1335 -338
rect 1503 -372 1515 -338
rect 1323 -378 1515 -372
rect 1581 -338 1773 -332
rect 1581 -372 1593 -338
rect 1761 -372 1773 -338
rect 1581 -378 1773 -372
rect 1839 -338 2031 -332
rect 1839 -372 1851 -338
rect 2019 -372 2031 -338
rect 1839 -378 2031 -372
rect 2097 -338 2289 -332
rect 2097 -372 2109 -338
rect 2277 -372 2289 -338
rect 2097 -378 2289 -372
rect 2355 -338 2547 -332
rect 2355 -372 2367 -338
rect 2535 -372 2547 -338
rect 2355 -378 2547 -372
<< properties >>
string FIXED_BBOX -2714 -493 2714 493
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
