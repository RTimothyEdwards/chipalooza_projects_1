* NGSPICE file created from isolated_switch.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6 w_n387_n462# a_29_n261# a_n129_n261# a_n29_n164#
+ a_n187_n164# a_129_n164#
X0 a_129_n164# a_29_n261# a_n29_n164# w_n387_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n164# a_n129_n261# a_n187_n164# w_n387_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HRGQF2 a_n321_n622# a_n29_n400# a_n187_n400#
+ a_129_n400# a_29_n488# a_n129_n488#
X0 a_n29_n400# a_n129_n488# a_n187_n400# a_n321_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_129_n400# a_29_n488# a_n29_n400# a_n321_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U62SY6 a_n187_n64# w_n387_n362# a_129_n64# a_29_n161#
+ a_n129_n161# a_n29_n64#
X0 a_129_n64# a_29_n161# a_n29_n64# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n64# a_n129_n161# a_n187_n64# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4 a_n242_n622# a_50_n400# a_n108_n400# a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n242_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6 a_n108_n164# a_n50_n261# w_n308_n462#
+ a_50_n164#
X0 a_50_n164# a_n50_n261# a_n108_n164# w_n308_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ3N a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RK a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt isolated_switch on vss out in vdd
Xsky130_fd_pr__pfet_g5v0d10v5_U6V9Y6_0 vdd onb onb m1_1166_n2330# out out sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6
Xsky130_fd_pr__nfet_g5v0d10v5_HRGQF2_0 vss m1_1166_n2330# out out onp onp sky130_fd_pr__nfet_g5v0d10v5_HRGQF2
Xsky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 onb vdd onb on on vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM1 vss in m1_1166_n2330# m1_1166_n2330# onp onp sky130_fd_pr__nfet_g5v0d10v5_HRGQF2
XXM3 vss in in onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
XXM4 vdd onb onb in m1_1166_n2330# m1_1166_n2330# sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6
XXM5 vss m1_1166_n2330# m1_1166_n2330# onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
XXM6 m1_1166_n2330# onp vdd m1_1166_n2330# sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
XXM7 onp vdd onp onb onb vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
Xsky130_fd_pr__nfet_g5v0d10v5_UNEQ3N_0 vss vss m1_1166_n2330# onb sky130_fd_pr__nfet_g5v0d10v5_UNEQ3N
XXM8 onp vss vss onb sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXD1 vss on sky130_fd_pr__diode_pw2nd_05v5_FT76RK
Xsky130_fd_pr__nfet_g5v0d10v5_MJGQJ4_0 vss m1_1166_n2330# m1_1166_n2330# onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
Xsky130_fd_pr__nfet_g5v0d10v5_MJGQJ4_1 vss out out onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
Xsky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_0 in onp vdd in sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
Xsky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_1 m1_1166_n2330# onp vdd m1_1166_n2330# sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
Xsky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_2 out onp vdd out sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
XXM10 onb vss vss on sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
.ends

