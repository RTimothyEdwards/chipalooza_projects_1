magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< error_p >>
rect -7017 1566 7017 1600
rect -7047 -1566 7047 1566
rect -7017 -1600 7017 -1566
<< nwell >>
rect -7017 -1600 7017 1600
<< mvpmos >>
rect -6923 -1500 -6823 1500
rect -6765 -1500 -6665 1500
rect -6607 -1500 -6507 1500
rect -6449 -1500 -6349 1500
rect -6291 -1500 -6191 1500
rect -6133 -1500 -6033 1500
rect -5975 -1500 -5875 1500
rect -5817 -1500 -5717 1500
rect -5659 -1500 -5559 1500
rect -5501 -1500 -5401 1500
rect -5343 -1500 -5243 1500
rect -5185 -1500 -5085 1500
rect -5027 -1500 -4927 1500
rect -4869 -1500 -4769 1500
rect -4711 -1500 -4611 1500
rect -4553 -1500 -4453 1500
rect -4395 -1500 -4295 1500
rect -4237 -1500 -4137 1500
rect -4079 -1500 -3979 1500
rect -3921 -1500 -3821 1500
rect -3763 -1500 -3663 1500
rect -3605 -1500 -3505 1500
rect -3447 -1500 -3347 1500
rect -3289 -1500 -3189 1500
rect -3131 -1500 -3031 1500
rect -2973 -1500 -2873 1500
rect -2815 -1500 -2715 1500
rect -2657 -1500 -2557 1500
rect -2499 -1500 -2399 1500
rect -2341 -1500 -2241 1500
rect -2183 -1500 -2083 1500
rect -2025 -1500 -1925 1500
rect -1867 -1500 -1767 1500
rect -1709 -1500 -1609 1500
rect -1551 -1500 -1451 1500
rect -1393 -1500 -1293 1500
rect -1235 -1500 -1135 1500
rect -1077 -1500 -977 1500
rect -919 -1500 -819 1500
rect -761 -1500 -661 1500
rect -603 -1500 -503 1500
rect -445 -1500 -345 1500
rect -287 -1500 -187 1500
rect -129 -1500 -29 1500
rect 29 -1500 129 1500
rect 187 -1500 287 1500
rect 345 -1500 445 1500
rect 503 -1500 603 1500
rect 661 -1500 761 1500
rect 819 -1500 919 1500
rect 977 -1500 1077 1500
rect 1135 -1500 1235 1500
rect 1293 -1500 1393 1500
rect 1451 -1500 1551 1500
rect 1609 -1500 1709 1500
rect 1767 -1500 1867 1500
rect 1925 -1500 2025 1500
rect 2083 -1500 2183 1500
rect 2241 -1500 2341 1500
rect 2399 -1500 2499 1500
rect 2557 -1500 2657 1500
rect 2715 -1500 2815 1500
rect 2873 -1500 2973 1500
rect 3031 -1500 3131 1500
rect 3189 -1500 3289 1500
rect 3347 -1500 3447 1500
rect 3505 -1500 3605 1500
rect 3663 -1500 3763 1500
rect 3821 -1500 3921 1500
rect 3979 -1500 4079 1500
rect 4137 -1500 4237 1500
rect 4295 -1500 4395 1500
rect 4453 -1500 4553 1500
rect 4611 -1500 4711 1500
rect 4769 -1500 4869 1500
rect 4927 -1500 5027 1500
rect 5085 -1500 5185 1500
rect 5243 -1500 5343 1500
rect 5401 -1500 5501 1500
rect 5559 -1500 5659 1500
rect 5717 -1500 5817 1500
rect 5875 -1500 5975 1500
rect 6033 -1500 6133 1500
rect 6191 -1500 6291 1500
rect 6349 -1500 6449 1500
rect 6507 -1500 6607 1500
rect 6665 -1500 6765 1500
rect 6823 -1500 6923 1500
<< mvpdiff >>
rect -6981 1488 -6923 1500
rect -6981 -1488 -6969 1488
rect -6935 -1488 -6923 1488
rect -6981 -1500 -6923 -1488
rect -6823 1488 -6765 1500
rect -6823 -1488 -6811 1488
rect -6777 -1488 -6765 1488
rect -6823 -1500 -6765 -1488
rect -6665 1488 -6607 1500
rect -6665 -1488 -6653 1488
rect -6619 -1488 -6607 1488
rect -6665 -1500 -6607 -1488
rect -6507 1488 -6449 1500
rect -6507 -1488 -6495 1488
rect -6461 -1488 -6449 1488
rect -6507 -1500 -6449 -1488
rect -6349 1488 -6291 1500
rect -6349 -1488 -6337 1488
rect -6303 -1488 -6291 1488
rect -6349 -1500 -6291 -1488
rect -6191 1488 -6133 1500
rect -6191 -1488 -6179 1488
rect -6145 -1488 -6133 1488
rect -6191 -1500 -6133 -1488
rect -6033 1488 -5975 1500
rect -6033 -1488 -6021 1488
rect -5987 -1488 -5975 1488
rect -6033 -1500 -5975 -1488
rect -5875 1488 -5817 1500
rect -5875 -1488 -5863 1488
rect -5829 -1488 -5817 1488
rect -5875 -1500 -5817 -1488
rect -5717 1488 -5659 1500
rect -5717 -1488 -5705 1488
rect -5671 -1488 -5659 1488
rect -5717 -1500 -5659 -1488
rect -5559 1488 -5501 1500
rect -5559 -1488 -5547 1488
rect -5513 -1488 -5501 1488
rect -5559 -1500 -5501 -1488
rect -5401 1488 -5343 1500
rect -5401 -1488 -5389 1488
rect -5355 -1488 -5343 1488
rect -5401 -1500 -5343 -1488
rect -5243 1488 -5185 1500
rect -5243 -1488 -5231 1488
rect -5197 -1488 -5185 1488
rect -5243 -1500 -5185 -1488
rect -5085 1488 -5027 1500
rect -5085 -1488 -5073 1488
rect -5039 -1488 -5027 1488
rect -5085 -1500 -5027 -1488
rect -4927 1488 -4869 1500
rect -4927 -1488 -4915 1488
rect -4881 -1488 -4869 1488
rect -4927 -1500 -4869 -1488
rect -4769 1488 -4711 1500
rect -4769 -1488 -4757 1488
rect -4723 -1488 -4711 1488
rect -4769 -1500 -4711 -1488
rect -4611 1488 -4553 1500
rect -4611 -1488 -4599 1488
rect -4565 -1488 -4553 1488
rect -4611 -1500 -4553 -1488
rect -4453 1488 -4395 1500
rect -4453 -1488 -4441 1488
rect -4407 -1488 -4395 1488
rect -4453 -1500 -4395 -1488
rect -4295 1488 -4237 1500
rect -4295 -1488 -4283 1488
rect -4249 -1488 -4237 1488
rect -4295 -1500 -4237 -1488
rect -4137 1488 -4079 1500
rect -4137 -1488 -4125 1488
rect -4091 -1488 -4079 1488
rect -4137 -1500 -4079 -1488
rect -3979 1488 -3921 1500
rect -3979 -1488 -3967 1488
rect -3933 -1488 -3921 1488
rect -3979 -1500 -3921 -1488
rect -3821 1488 -3763 1500
rect -3821 -1488 -3809 1488
rect -3775 -1488 -3763 1488
rect -3821 -1500 -3763 -1488
rect -3663 1488 -3605 1500
rect -3663 -1488 -3651 1488
rect -3617 -1488 -3605 1488
rect -3663 -1500 -3605 -1488
rect -3505 1488 -3447 1500
rect -3505 -1488 -3493 1488
rect -3459 -1488 -3447 1488
rect -3505 -1500 -3447 -1488
rect -3347 1488 -3289 1500
rect -3347 -1488 -3335 1488
rect -3301 -1488 -3289 1488
rect -3347 -1500 -3289 -1488
rect -3189 1488 -3131 1500
rect -3189 -1488 -3177 1488
rect -3143 -1488 -3131 1488
rect -3189 -1500 -3131 -1488
rect -3031 1488 -2973 1500
rect -3031 -1488 -3019 1488
rect -2985 -1488 -2973 1488
rect -3031 -1500 -2973 -1488
rect -2873 1488 -2815 1500
rect -2873 -1488 -2861 1488
rect -2827 -1488 -2815 1488
rect -2873 -1500 -2815 -1488
rect -2715 1488 -2657 1500
rect -2715 -1488 -2703 1488
rect -2669 -1488 -2657 1488
rect -2715 -1500 -2657 -1488
rect -2557 1488 -2499 1500
rect -2557 -1488 -2545 1488
rect -2511 -1488 -2499 1488
rect -2557 -1500 -2499 -1488
rect -2399 1488 -2341 1500
rect -2399 -1488 -2387 1488
rect -2353 -1488 -2341 1488
rect -2399 -1500 -2341 -1488
rect -2241 1488 -2183 1500
rect -2241 -1488 -2229 1488
rect -2195 -1488 -2183 1488
rect -2241 -1500 -2183 -1488
rect -2083 1488 -2025 1500
rect -2083 -1488 -2071 1488
rect -2037 -1488 -2025 1488
rect -2083 -1500 -2025 -1488
rect -1925 1488 -1867 1500
rect -1925 -1488 -1913 1488
rect -1879 -1488 -1867 1488
rect -1925 -1500 -1867 -1488
rect -1767 1488 -1709 1500
rect -1767 -1488 -1755 1488
rect -1721 -1488 -1709 1488
rect -1767 -1500 -1709 -1488
rect -1609 1488 -1551 1500
rect -1609 -1488 -1597 1488
rect -1563 -1488 -1551 1488
rect -1609 -1500 -1551 -1488
rect -1451 1488 -1393 1500
rect -1451 -1488 -1439 1488
rect -1405 -1488 -1393 1488
rect -1451 -1500 -1393 -1488
rect -1293 1488 -1235 1500
rect -1293 -1488 -1281 1488
rect -1247 -1488 -1235 1488
rect -1293 -1500 -1235 -1488
rect -1135 1488 -1077 1500
rect -1135 -1488 -1123 1488
rect -1089 -1488 -1077 1488
rect -1135 -1500 -1077 -1488
rect -977 1488 -919 1500
rect -977 -1488 -965 1488
rect -931 -1488 -919 1488
rect -977 -1500 -919 -1488
rect -819 1488 -761 1500
rect -819 -1488 -807 1488
rect -773 -1488 -761 1488
rect -819 -1500 -761 -1488
rect -661 1488 -603 1500
rect -661 -1488 -649 1488
rect -615 -1488 -603 1488
rect -661 -1500 -603 -1488
rect -503 1488 -445 1500
rect -503 -1488 -491 1488
rect -457 -1488 -445 1488
rect -503 -1500 -445 -1488
rect -345 1488 -287 1500
rect -345 -1488 -333 1488
rect -299 -1488 -287 1488
rect -345 -1500 -287 -1488
rect -187 1488 -129 1500
rect -187 -1488 -175 1488
rect -141 -1488 -129 1488
rect -187 -1500 -129 -1488
rect -29 1488 29 1500
rect -29 -1488 -17 1488
rect 17 -1488 29 1488
rect -29 -1500 29 -1488
rect 129 1488 187 1500
rect 129 -1488 141 1488
rect 175 -1488 187 1488
rect 129 -1500 187 -1488
rect 287 1488 345 1500
rect 287 -1488 299 1488
rect 333 -1488 345 1488
rect 287 -1500 345 -1488
rect 445 1488 503 1500
rect 445 -1488 457 1488
rect 491 -1488 503 1488
rect 445 -1500 503 -1488
rect 603 1488 661 1500
rect 603 -1488 615 1488
rect 649 -1488 661 1488
rect 603 -1500 661 -1488
rect 761 1488 819 1500
rect 761 -1488 773 1488
rect 807 -1488 819 1488
rect 761 -1500 819 -1488
rect 919 1488 977 1500
rect 919 -1488 931 1488
rect 965 -1488 977 1488
rect 919 -1500 977 -1488
rect 1077 1488 1135 1500
rect 1077 -1488 1089 1488
rect 1123 -1488 1135 1488
rect 1077 -1500 1135 -1488
rect 1235 1488 1293 1500
rect 1235 -1488 1247 1488
rect 1281 -1488 1293 1488
rect 1235 -1500 1293 -1488
rect 1393 1488 1451 1500
rect 1393 -1488 1405 1488
rect 1439 -1488 1451 1488
rect 1393 -1500 1451 -1488
rect 1551 1488 1609 1500
rect 1551 -1488 1563 1488
rect 1597 -1488 1609 1488
rect 1551 -1500 1609 -1488
rect 1709 1488 1767 1500
rect 1709 -1488 1721 1488
rect 1755 -1488 1767 1488
rect 1709 -1500 1767 -1488
rect 1867 1488 1925 1500
rect 1867 -1488 1879 1488
rect 1913 -1488 1925 1488
rect 1867 -1500 1925 -1488
rect 2025 1488 2083 1500
rect 2025 -1488 2037 1488
rect 2071 -1488 2083 1488
rect 2025 -1500 2083 -1488
rect 2183 1488 2241 1500
rect 2183 -1488 2195 1488
rect 2229 -1488 2241 1488
rect 2183 -1500 2241 -1488
rect 2341 1488 2399 1500
rect 2341 -1488 2353 1488
rect 2387 -1488 2399 1488
rect 2341 -1500 2399 -1488
rect 2499 1488 2557 1500
rect 2499 -1488 2511 1488
rect 2545 -1488 2557 1488
rect 2499 -1500 2557 -1488
rect 2657 1488 2715 1500
rect 2657 -1488 2669 1488
rect 2703 -1488 2715 1488
rect 2657 -1500 2715 -1488
rect 2815 1488 2873 1500
rect 2815 -1488 2827 1488
rect 2861 -1488 2873 1488
rect 2815 -1500 2873 -1488
rect 2973 1488 3031 1500
rect 2973 -1488 2985 1488
rect 3019 -1488 3031 1488
rect 2973 -1500 3031 -1488
rect 3131 1488 3189 1500
rect 3131 -1488 3143 1488
rect 3177 -1488 3189 1488
rect 3131 -1500 3189 -1488
rect 3289 1488 3347 1500
rect 3289 -1488 3301 1488
rect 3335 -1488 3347 1488
rect 3289 -1500 3347 -1488
rect 3447 1488 3505 1500
rect 3447 -1488 3459 1488
rect 3493 -1488 3505 1488
rect 3447 -1500 3505 -1488
rect 3605 1488 3663 1500
rect 3605 -1488 3617 1488
rect 3651 -1488 3663 1488
rect 3605 -1500 3663 -1488
rect 3763 1488 3821 1500
rect 3763 -1488 3775 1488
rect 3809 -1488 3821 1488
rect 3763 -1500 3821 -1488
rect 3921 1488 3979 1500
rect 3921 -1488 3933 1488
rect 3967 -1488 3979 1488
rect 3921 -1500 3979 -1488
rect 4079 1488 4137 1500
rect 4079 -1488 4091 1488
rect 4125 -1488 4137 1488
rect 4079 -1500 4137 -1488
rect 4237 1488 4295 1500
rect 4237 -1488 4249 1488
rect 4283 -1488 4295 1488
rect 4237 -1500 4295 -1488
rect 4395 1488 4453 1500
rect 4395 -1488 4407 1488
rect 4441 -1488 4453 1488
rect 4395 -1500 4453 -1488
rect 4553 1488 4611 1500
rect 4553 -1488 4565 1488
rect 4599 -1488 4611 1488
rect 4553 -1500 4611 -1488
rect 4711 1488 4769 1500
rect 4711 -1488 4723 1488
rect 4757 -1488 4769 1488
rect 4711 -1500 4769 -1488
rect 4869 1488 4927 1500
rect 4869 -1488 4881 1488
rect 4915 -1488 4927 1488
rect 4869 -1500 4927 -1488
rect 5027 1488 5085 1500
rect 5027 -1488 5039 1488
rect 5073 -1488 5085 1488
rect 5027 -1500 5085 -1488
rect 5185 1488 5243 1500
rect 5185 -1488 5197 1488
rect 5231 -1488 5243 1488
rect 5185 -1500 5243 -1488
rect 5343 1488 5401 1500
rect 5343 -1488 5355 1488
rect 5389 -1488 5401 1488
rect 5343 -1500 5401 -1488
rect 5501 1488 5559 1500
rect 5501 -1488 5513 1488
rect 5547 -1488 5559 1488
rect 5501 -1500 5559 -1488
rect 5659 1488 5717 1500
rect 5659 -1488 5671 1488
rect 5705 -1488 5717 1488
rect 5659 -1500 5717 -1488
rect 5817 1488 5875 1500
rect 5817 -1488 5829 1488
rect 5863 -1488 5875 1488
rect 5817 -1500 5875 -1488
rect 5975 1488 6033 1500
rect 5975 -1488 5987 1488
rect 6021 -1488 6033 1488
rect 5975 -1500 6033 -1488
rect 6133 1488 6191 1500
rect 6133 -1488 6145 1488
rect 6179 -1488 6191 1488
rect 6133 -1500 6191 -1488
rect 6291 1488 6349 1500
rect 6291 -1488 6303 1488
rect 6337 -1488 6349 1488
rect 6291 -1500 6349 -1488
rect 6449 1488 6507 1500
rect 6449 -1488 6461 1488
rect 6495 -1488 6507 1488
rect 6449 -1500 6507 -1488
rect 6607 1488 6665 1500
rect 6607 -1488 6619 1488
rect 6653 -1488 6665 1488
rect 6607 -1500 6665 -1488
rect 6765 1488 6823 1500
rect 6765 -1488 6777 1488
rect 6811 -1488 6823 1488
rect 6765 -1500 6823 -1488
rect 6923 1488 6981 1500
rect 6923 -1488 6935 1488
rect 6969 -1488 6981 1488
rect 6923 -1500 6981 -1488
<< mvpdiffc >>
rect -6969 -1488 -6935 1488
rect -6811 -1488 -6777 1488
rect -6653 -1488 -6619 1488
rect -6495 -1488 -6461 1488
rect -6337 -1488 -6303 1488
rect -6179 -1488 -6145 1488
rect -6021 -1488 -5987 1488
rect -5863 -1488 -5829 1488
rect -5705 -1488 -5671 1488
rect -5547 -1488 -5513 1488
rect -5389 -1488 -5355 1488
rect -5231 -1488 -5197 1488
rect -5073 -1488 -5039 1488
rect -4915 -1488 -4881 1488
rect -4757 -1488 -4723 1488
rect -4599 -1488 -4565 1488
rect -4441 -1488 -4407 1488
rect -4283 -1488 -4249 1488
rect -4125 -1488 -4091 1488
rect -3967 -1488 -3933 1488
rect -3809 -1488 -3775 1488
rect -3651 -1488 -3617 1488
rect -3493 -1488 -3459 1488
rect -3335 -1488 -3301 1488
rect -3177 -1488 -3143 1488
rect -3019 -1488 -2985 1488
rect -2861 -1488 -2827 1488
rect -2703 -1488 -2669 1488
rect -2545 -1488 -2511 1488
rect -2387 -1488 -2353 1488
rect -2229 -1488 -2195 1488
rect -2071 -1488 -2037 1488
rect -1913 -1488 -1879 1488
rect -1755 -1488 -1721 1488
rect -1597 -1488 -1563 1488
rect -1439 -1488 -1405 1488
rect -1281 -1488 -1247 1488
rect -1123 -1488 -1089 1488
rect -965 -1488 -931 1488
rect -807 -1488 -773 1488
rect -649 -1488 -615 1488
rect -491 -1488 -457 1488
rect -333 -1488 -299 1488
rect -175 -1488 -141 1488
rect -17 -1488 17 1488
rect 141 -1488 175 1488
rect 299 -1488 333 1488
rect 457 -1488 491 1488
rect 615 -1488 649 1488
rect 773 -1488 807 1488
rect 931 -1488 965 1488
rect 1089 -1488 1123 1488
rect 1247 -1488 1281 1488
rect 1405 -1488 1439 1488
rect 1563 -1488 1597 1488
rect 1721 -1488 1755 1488
rect 1879 -1488 1913 1488
rect 2037 -1488 2071 1488
rect 2195 -1488 2229 1488
rect 2353 -1488 2387 1488
rect 2511 -1488 2545 1488
rect 2669 -1488 2703 1488
rect 2827 -1488 2861 1488
rect 2985 -1488 3019 1488
rect 3143 -1488 3177 1488
rect 3301 -1488 3335 1488
rect 3459 -1488 3493 1488
rect 3617 -1488 3651 1488
rect 3775 -1488 3809 1488
rect 3933 -1488 3967 1488
rect 4091 -1488 4125 1488
rect 4249 -1488 4283 1488
rect 4407 -1488 4441 1488
rect 4565 -1488 4599 1488
rect 4723 -1488 4757 1488
rect 4881 -1488 4915 1488
rect 5039 -1488 5073 1488
rect 5197 -1488 5231 1488
rect 5355 -1488 5389 1488
rect 5513 -1488 5547 1488
rect 5671 -1488 5705 1488
rect 5829 -1488 5863 1488
rect 5987 -1488 6021 1488
rect 6145 -1488 6179 1488
rect 6303 -1488 6337 1488
rect 6461 -1488 6495 1488
rect 6619 -1488 6653 1488
rect 6777 -1488 6811 1488
rect 6935 -1488 6969 1488
<< poly >>
rect -6923 1581 -6823 1597
rect -6923 1547 -6907 1581
rect -6839 1547 -6823 1581
rect -6923 1500 -6823 1547
rect -6765 1581 -6665 1597
rect -6765 1547 -6749 1581
rect -6681 1547 -6665 1581
rect -6765 1500 -6665 1547
rect -6607 1581 -6507 1597
rect -6607 1547 -6591 1581
rect -6523 1547 -6507 1581
rect -6607 1500 -6507 1547
rect -6449 1581 -6349 1597
rect -6449 1547 -6433 1581
rect -6365 1547 -6349 1581
rect -6449 1500 -6349 1547
rect -6291 1581 -6191 1597
rect -6291 1547 -6275 1581
rect -6207 1547 -6191 1581
rect -6291 1500 -6191 1547
rect -6133 1581 -6033 1597
rect -6133 1547 -6117 1581
rect -6049 1547 -6033 1581
rect -6133 1500 -6033 1547
rect -5975 1581 -5875 1597
rect -5975 1547 -5959 1581
rect -5891 1547 -5875 1581
rect -5975 1500 -5875 1547
rect -5817 1581 -5717 1597
rect -5817 1547 -5801 1581
rect -5733 1547 -5717 1581
rect -5817 1500 -5717 1547
rect -5659 1581 -5559 1597
rect -5659 1547 -5643 1581
rect -5575 1547 -5559 1581
rect -5659 1500 -5559 1547
rect -5501 1581 -5401 1597
rect -5501 1547 -5485 1581
rect -5417 1547 -5401 1581
rect -5501 1500 -5401 1547
rect -5343 1581 -5243 1597
rect -5343 1547 -5327 1581
rect -5259 1547 -5243 1581
rect -5343 1500 -5243 1547
rect -5185 1581 -5085 1597
rect -5185 1547 -5169 1581
rect -5101 1547 -5085 1581
rect -5185 1500 -5085 1547
rect -5027 1581 -4927 1597
rect -5027 1547 -5011 1581
rect -4943 1547 -4927 1581
rect -5027 1500 -4927 1547
rect -4869 1581 -4769 1597
rect -4869 1547 -4853 1581
rect -4785 1547 -4769 1581
rect -4869 1500 -4769 1547
rect -4711 1581 -4611 1597
rect -4711 1547 -4695 1581
rect -4627 1547 -4611 1581
rect -4711 1500 -4611 1547
rect -4553 1581 -4453 1597
rect -4553 1547 -4537 1581
rect -4469 1547 -4453 1581
rect -4553 1500 -4453 1547
rect -4395 1581 -4295 1597
rect -4395 1547 -4379 1581
rect -4311 1547 -4295 1581
rect -4395 1500 -4295 1547
rect -4237 1581 -4137 1597
rect -4237 1547 -4221 1581
rect -4153 1547 -4137 1581
rect -4237 1500 -4137 1547
rect -4079 1581 -3979 1597
rect -4079 1547 -4063 1581
rect -3995 1547 -3979 1581
rect -4079 1500 -3979 1547
rect -3921 1581 -3821 1597
rect -3921 1547 -3905 1581
rect -3837 1547 -3821 1581
rect -3921 1500 -3821 1547
rect -3763 1581 -3663 1597
rect -3763 1547 -3747 1581
rect -3679 1547 -3663 1581
rect -3763 1500 -3663 1547
rect -3605 1581 -3505 1597
rect -3605 1547 -3589 1581
rect -3521 1547 -3505 1581
rect -3605 1500 -3505 1547
rect -3447 1581 -3347 1597
rect -3447 1547 -3431 1581
rect -3363 1547 -3347 1581
rect -3447 1500 -3347 1547
rect -3289 1581 -3189 1597
rect -3289 1547 -3273 1581
rect -3205 1547 -3189 1581
rect -3289 1500 -3189 1547
rect -3131 1581 -3031 1597
rect -3131 1547 -3115 1581
rect -3047 1547 -3031 1581
rect -3131 1500 -3031 1547
rect -2973 1581 -2873 1597
rect -2973 1547 -2957 1581
rect -2889 1547 -2873 1581
rect -2973 1500 -2873 1547
rect -2815 1581 -2715 1597
rect -2815 1547 -2799 1581
rect -2731 1547 -2715 1581
rect -2815 1500 -2715 1547
rect -2657 1581 -2557 1597
rect -2657 1547 -2641 1581
rect -2573 1547 -2557 1581
rect -2657 1500 -2557 1547
rect -2499 1581 -2399 1597
rect -2499 1547 -2483 1581
rect -2415 1547 -2399 1581
rect -2499 1500 -2399 1547
rect -2341 1581 -2241 1597
rect -2341 1547 -2325 1581
rect -2257 1547 -2241 1581
rect -2341 1500 -2241 1547
rect -2183 1581 -2083 1597
rect -2183 1547 -2167 1581
rect -2099 1547 -2083 1581
rect -2183 1500 -2083 1547
rect -2025 1581 -1925 1597
rect -2025 1547 -2009 1581
rect -1941 1547 -1925 1581
rect -2025 1500 -1925 1547
rect -1867 1581 -1767 1597
rect -1867 1547 -1851 1581
rect -1783 1547 -1767 1581
rect -1867 1500 -1767 1547
rect -1709 1581 -1609 1597
rect -1709 1547 -1693 1581
rect -1625 1547 -1609 1581
rect -1709 1500 -1609 1547
rect -1551 1581 -1451 1597
rect -1551 1547 -1535 1581
rect -1467 1547 -1451 1581
rect -1551 1500 -1451 1547
rect -1393 1581 -1293 1597
rect -1393 1547 -1377 1581
rect -1309 1547 -1293 1581
rect -1393 1500 -1293 1547
rect -1235 1581 -1135 1597
rect -1235 1547 -1219 1581
rect -1151 1547 -1135 1581
rect -1235 1500 -1135 1547
rect -1077 1581 -977 1597
rect -1077 1547 -1061 1581
rect -993 1547 -977 1581
rect -1077 1500 -977 1547
rect -919 1581 -819 1597
rect -919 1547 -903 1581
rect -835 1547 -819 1581
rect -919 1500 -819 1547
rect -761 1581 -661 1597
rect -761 1547 -745 1581
rect -677 1547 -661 1581
rect -761 1500 -661 1547
rect -603 1581 -503 1597
rect -603 1547 -587 1581
rect -519 1547 -503 1581
rect -603 1500 -503 1547
rect -445 1581 -345 1597
rect -445 1547 -429 1581
rect -361 1547 -345 1581
rect -445 1500 -345 1547
rect -287 1581 -187 1597
rect -287 1547 -271 1581
rect -203 1547 -187 1581
rect -287 1500 -187 1547
rect -129 1581 -29 1597
rect -129 1547 -113 1581
rect -45 1547 -29 1581
rect -129 1500 -29 1547
rect 29 1581 129 1597
rect 29 1547 45 1581
rect 113 1547 129 1581
rect 29 1500 129 1547
rect 187 1581 287 1597
rect 187 1547 203 1581
rect 271 1547 287 1581
rect 187 1500 287 1547
rect 345 1581 445 1597
rect 345 1547 361 1581
rect 429 1547 445 1581
rect 345 1500 445 1547
rect 503 1581 603 1597
rect 503 1547 519 1581
rect 587 1547 603 1581
rect 503 1500 603 1547
rect 661 1581 761 1597
rect 661 1547 677 1581
rect 745 1547 761 1581
rect 661 1500 761 1547
rect 819 1581 919 1597
rect 819 1547 835 1581
rect 903 1547 919 1581
rect 819 1500 919 1547
rect 977 1581 1077 1597
rect 977 1547 993 1581
rect 1061 1547 1077 1581
rect 977 1500 1077 1547
rect 1135 1581 1235 1597
rect 1135 1547 1151 1581
rect 1219 1547 1235 1581
rect 1135 1500 1235 1547
rect 1293 1581 1393 1597
rect 1293 1547 1309 1581
rect 1377 1547 1393 1581
rect 1293 1500 1393 1547
rect 1451 1581 1551 1597
rect 1451 1547 1467 1581
rect 1535 1547 1551 1581
rect 1451 1500 1551 1547
rect 1609 1581 1709 1597
rect 1609 1547 1625 1581
rect 1693 1547 1709 1581
rect 1609 1500 1709 1547
rect 1767 1581 1867 1597
rect 1767 1547 1783 1581
rect 1851 1547 1867 1581
rect 1767 1500 1867 1547
rect 1925 1581 2025 1597
rect 1925 1547 1941 1581
rect 2009 1547 2025 1581
rect 1925 1500 2025 1547
rect 2083 1581 2183 1597
rect 2083 1547 2099 1581
rect 2167 1547 2183 1581
rect 2083 1500 2183 1547
rect 2241 1581 2341 1597
rect 2241 1547 2257 1581
rect 2325 1547 2341 1581
rect 2241 1500 2341 1547
rect 2399 1581 2499 1597
rect 2399 1547 2415 1581
rect 2483 1547 2499 1581
rect 2399 1500 2499 1547
rect 2557 1581 2657 1597
rect 2557 1547 2573 1581
rect 2641 1547 2657 1581
rect 2557 1500 2657 1547
rect 2715 1581 2815 1597
rect 2715 1547 2731 1581
rect 2799 1547 2815 1581
rect 2715 1500 2815 1547
rect 2873 1581 2973 1597
rect 2873 1547 2889 1581
rect 2957 1547 2973 1581
rect 2873 1500 2973 1547
rect 3031 1581 3131 1597
rect 3031 1547 3047 1581
rect 3115 1547 3131 1581
rect 3031 1500 3131 1547
rect 3189 1581 3289 1597
rect 3189 1547 3205 1581
rect 3273 1547 3289 1581
rect 3189 1500 3289 1547
rect 3347 1581 3447 1597
rect 3347 1547 3363 1581
rect 3431 1547 3447 1581
rect 3347 1500 3447 1547
rect 3505 1581 3605 1597
rect 3505 1547 3521 1581
rect 3589 1547 3605 1581
rect 3505 1500 3605 1547
rect 3663 1581 3763 1597
rect 3663 1547 3679 1581
rect 3747 1547 3763 1581
rect 3663 1500 3763 1547
rect 3821 1581 3921 1597
rect 3821 1547 3837 1581
rect 3905 1547 3921 1581
rect 3821 1500 3921 1547
rect 3979 1581 4079 1597
rect 3979 1547 3995 1581
rect 4063 1547 4079 1581
rect 3979 1500 4079 1547
rect 4137 1581 4237 1597
rect 4137 1547 4153 1581
rect 4221 1547 4237 1581
rect 4137 1500 4237 1547
rect 4295 1581 4395 1597
rect 4295 1547 4311 1581
rect 4379 1547 4395 1581
rect 4295 1500 4395 1547
rect 4453 1581 4553 1597
rect 4453 1547 4469 1581
rect 4537 1547 4553 1581
rect 4453 1500 4553 1547
rect 4611 1581 4711 1597
rect 4611 1547 4627 1581
rect 4695 1547 4711 1581
rect 4611 1500 4711 1547
rect 4769 1581 4869 1597
rect 4769 1547 4785 1581
rect 4853 1547 4869 1581
rect 4769 1500 4869 1547
rect 4927 1581 5027 1597
rect 4927 1547 4943 1581
rect 5011 1547 5027 1581
rect 4927 1500 5027 1547
rect 5085 1581 5185 1597
rect 5085 1547 5101 1581
rect 5169 1547 5185 1581
rect 5085 1500 5185 1547
rect 5243 1581 5343 1597
rect 5243 1547 5259 1581
rect 5327 1547 5343 1581
rect 5243 1500 5343 1547
rect 5401 1581 5501 1597
rect 5401 1547 5417 1581
rect 5485 1547 5501 1581
rect 5401 1500 5501 1547
rect 5559 1581 5659 1597
rect 5559 1547 5575 1581
rect 5643 1547 5659 1581
rect 5559 1500 5659 1547
rect 5717 1581 5817 1597
rect 5717 1547 5733 1581
rect 5801 1547 5817 1581
rect 5717 1500 5817 1547
rect 5875 1581 5975 1597
rect 5875 1547 5891 1581
rect 5959 1547 5975 1581
rect 5875 1500 5975 1547
rect 6033 1581 6133 1597
rect 6033 1547 6049 1581
rect 6117 1547 6133 1581
rect 6033 1500 6133 1547
rect 6191 1581 6291 1597
rect 6191 1547 6207 1581
rect 6275 1547 6291 1581
rect 6191 1500 6291 1547
rect 6349 1581 6449 1597
rect 6349 1547 6365 1581
rect 6433 1547 6449 1581
rect 6349 1500 6449 1547
rect 6507 1581 6607 1597
rect 6507 1547 6523 1581
rect 6591 1547 6607 1581
rect 6507 1500 6607 1547
rect 6665 1581 6765 1597
rect 6665 1547 6681 1581
rect 6749 1547 6765 1581
rect 6665 1500 6765 1547
rect 6823 1581 6923 1597
rect 6823 1547 6839 1581
rect 6907 1547 6923 1581
rect 6823 1500 6923 1547
rect -6923 -1547 -6823 -1500
rect -6923 -1581 -6907 -1547
rect -6839 -1581 -6823 -1547
rect -6923 -1597 -6823 -1581
rect -6765 -1547 -6665 -1500
rect -6765 -1581 -6749 -1547
rect -6681 -1581 -6665 -1547
rect -6765 -1597 -6665 -1581
rect -6607 -1547 -6507 -1500
rect -6607 -1581 -6591 -1547
rect -6523 -1581 -6507 -1547
rect -6607 -1597 -6507 -1581
rect -6449 -1547 -6349 -1500
rect -6449 -1581 -6433 -1547
rect -6365 -1581 -6349 -1547
rect -6449 -1597 -6349 -1581
rect -6291 -1547 -6191 -1500
rect -6291 -1581 -6275 -1547
rect -6207 -1581 -6191 -1547
rect -6291 -1597 -6191 -1581
rect -6133 -1547 -6033 -1500
rect -6133 -1581 -6117 -1547
rect -6049 -1581 -6033 -1547
rect -6133 -1597 -6033 -1581
rect -5975 -1547 -5875 -1500
rect -5975 -1581 -5959 -1547
rect -5891 -1581 -5875 -1547
rect -5975 -1597 -5875 -1581
rect -5817 -1547 -5717 -1500
rect -5817 -1581 -5801 -1547
rect -5733 -1581 -5717 -1547
rect -5817 -1597 -5717 -1581
rect -5659 -1547 -5559 -1500
rect -5659 -1581 -5643 -1547
rect -5575 -1581 -5559 -1547
rect -5659 -1597 -5559 -1581
rect -5501 -1547 -5401 -1500
rect -5501 -1581 -5485 -1547
rect -5417 -1581 -5401 -1547
rect -5501 -1597 -5401 -1581
rect -5343 -1547 -5243 -1500
rect -5343 -1581 -5327 -1547
rect -5259 -1581 -5243 -1547
rect -5343 -1597 -5243 -1581
rect -5185 -1547 -5085 -1500
rect -5185 -1581 -5169 -1547
rect -5101 -1581 -5085 -1547
rect -5185 -1597 -5085 -1581
rect -5027 -1547 -4927 -1500
rect -5027 -1581 -5011 -1547
rect -4943 -1581 -4927 -1547
rect -5027 -1597 -4927 -1581
rect -4869 -1547 -4769 -1500
rect -4869 -1581 -4853 -1547
rect -4785 -1581 -4769 -1547
rect -4869 -1597 -4769 -1581
rect -4711 -1547 -4611 -1500
rect -4711 -1581 -4695 -1547
rect -4627 -1581 -4611 -1547
rect -4711 -1597 -4611 -1581
rect -4553 -1547 -4453 -1500
rect -4553 -1581 -4537 -1547
rect -4469 -1581 -4453 -1547
rect -4553 -1597 -4453 -1581
rect -4395 -1547 -4295 -1500
rect -4395 -1581 -4379 -1547
rect -4311 -1581 -4295 -1547
rect -4395 -1597 -4295 -1581
rect -4237 -1547 -4137 -1500
rect -4237 -1581 -4221 -1547
rect -4153 -1581 -4137 -1547
rect -4237 -1597 -4137 -1581
rect -4079 -1547 -3979 -1500
rect -4079 -1581 -4063 -1547
rect -3995 -1581 -3979 -1547
rect -4079 -1597 -3979 -1581
rect -3921 -1547 -3821 -1500
rect -3921 -1581 -3905 -1547
rect -3837 -1581 -3821 -1547
rect -3921 -1597 -3821 -1581
rect -3763 -1547 -3663 -1500
rect -3763 -1581 -3747 -1547
rect -3679 -1581 -3663 -1547
rect -3763 -1597 -3663 -1581
rect -3605 -1547 -3505 -1500
rect -3605 -1581 -3589 -1547
rect -3521 -1581 -3505 -1547
rect -3605 -1597 -3505 -1581
rect -3447 -1547 -3347 -1500
rect -3447 -1581 -3431 -1547
rect -3363 -1581 -3347 -1547
rect -3447 -1597 -3347 -1581
rect -3289 -1547 -3189 -1500
rect -3289 -1581 -3273 -1547
rect -3205 -1581 -3189 -1547
rect -3289 -1597 -3189 -1581
rect -3131 -1547 -3031 -1500
rect -3131 -1581 -3115 -1547
rect -3047 -1581 -3031 -1547
rect -3131 -1597 -3031 -1581
rect -2973 -1547 -2873 -1500
rect -2973 -1581 -2957 -1547
rect -2889 -1581 -2873 -1547
rect -2973 -1597 -2873 -1581
rect -2815 -1547 -2715 -1500
rect -2815 -1581 -2799 -1547
rect -2731 -1581 -2715 -1547
rect -2815 -1597 -2715 -1581
rect -2657 -1547 -2557 -1500
rect -2657 -1581 -2641 -1547
rect -2573 -1581 -2557 -1547
rect -2657 -1597 -2557 -1581
rect -2499 -1547 -2399 -1500
rect -2499 -1581 -2483 -1547
rect -2415 -1581 -2399 -1547
rect -2499 -1597 -2399 -1581
rect -2341 -1547 -2241 -1500
rect -2341 -1581 -2325 -1547
rect -2257 -1581 -2241 -1547
rect -2341 -1597 -2241 -1581
rect -2183 -1547 -2083 -1500
rect -2183 -1581 -2167 -1547
rect -2099 -1581 -2083 -1547
rect -2183 -1597 -2083 -1581
rect -2025 -1547 -1925 -1500
rect -2025 -1581 -2009 -1547
rect -1941 -1581 -1925 -1547
rect -2025 -1597 -1925 -1581
rect -1867 -1547 -1767 -1500
rect -1867 -1581 -1851 -1547
rect -1783 -1581 -1767 -1547
rect -1867 -1597 -1767 -1581
rect -1709 -1547 -1609 -1500
rect -1709 -1581 -1693 -1547
rect -1625 -1581 -1609 -1547
rect -1709 -1597 -1609 -1581
rect -1551 -1547 -1451 -1500
rect -1551 -1581 -1535 -1547
rect -1467 -1581 -1451 -1547
rect -1551 -1597 -1451 -1581
rect -1393 -1547 -1293 -1500
rect -1393 -1581 -1377 -1547
rect -1309 -1581 -1293 -1547
rect -1393 -1597 -1293 -1581
rect -1235 -1547 -1135 -1500
rect -1235 -1581 -1219 -1547
rect -1151 -1581 -1135 -1547
rect -1235 -1597 -1135 -1581
rect -1077 -1547 -977 -1500
rect -1077 -1581 -1061 -1547
rect -993 -1581 -977 -1547
rect -1077 -1597 -977 -1581
rect -919 -1547 -819 -1500
rect -919 -1581 -903 -1547
rect -835 -1581 -819 -1547
rect -919 -1597 -819 -1581
rect -761 -1547 -661 -1500
rect -761 -1581 -745 -1547
rect -677 -1581 -661 -1547
rect -761 -1597 -661 -1581
rect -603 -1547 -503 -1500
rect -603 -1581 -587 -1547
rect -519 -1581 -503 -1547
rect -603 -1597 -503 -1581
rect -445 -1547 -345 -1500
rect -445 -1581 -429 -1547
rect -361 -1581 -345 -1547
rect -445 -1597 -345 -1581
rect -287 -1547 -187 -1500
rect -287 -1581 -271 -1547
rect -203 -1581 -187 -1547
rect -287 -1597 -187 -1581
rect -129 -1547 -29 -1500
rect -129 -1581 -113 -1547
rect -45 -1581 -29 -1547
rect -129 -1597 -29 -1581
rect 29 -1547 129 -1500
rect 29 -1581 45 -1547
rect 113 -1581 129 -1547
rect 29 -1597 129 -1581
rect 187 -1547 287 -1500
rect 187 -1581 203 -1547
rect 271 -1581 287 -1547
rect 187 -1597 287 -1581
rect 345 -1547 445 -1500
rect 345 -1581 361 -1547
rect 429 -1581 445 -1547
rect 345 -1597 445 -1581
rect 503 -1547 603 -1500
rect 503 -1581 519 -1547
rect 587 -1581 603 -1547
rect 503 -1597 603 -1581
rect 661 -1547 761 -1500
rect 661 -1581 677 -1547
rect 745 -1581 761 -1547
rect 661 -1597 761 -1581
rect 819 -1547 919 -1500
rect 819 -1581 835 -1547
rect 903 -1581 919 -1547
rect 819 -1597 919 -1581
rect 977 -1547 1077 -1500
rect 977 -1581 993 -1547
rect 1061 -1581 1077 -1547
rect 977 -1597 1077 -1581
rect 1135 -1547 1235 -1500
rect 1135 -1581 1151 -1547
rect 1219 -1581 1235 -1547
rect 1135 -1597 1235 -1581
rect 1293 -1547 1393 -1500
rect 1293 -1581 1309 -1547
rect 1377 -1581 1393 -1547
rect 1293 -1597 1393 -1581
rect 1451 -1547 1551 -1500
rect 1451 -1581 1467 -1547
rect 1535 -1581 1551 -1547
rect 1451 -1597 1551 -1581
rect 1609 -1547 1709 -1500
rect 1609 -1581 1625 -1547
rect 1693 -1581 1709 -1547
rect 1609 -1597 1709 -1581
rect 1767 -1547 1867 -1500
rect 1767 -1581 1783 -1547
rect 1851 -1581 1867 -1547
rect 1767 -1597 1867 -1581
rect 1925 -1547 2025 -1500
rect 1925 -1581 1941 -1547
rect 2009 -1581 2025 -1547
rect 1925 -1597 2025 -1581
rect 2083 -1547 2183 -1500
rect 2083 -1581 2099 -1547
rect 2167 -1581 2183 -1547
rect 2083 -1597 2183 -1581
rect 2241 -1547 2341 -1500
rect 2241 -1581 2257 -1547
rect 2325 -1581 2341 -1547
rect 2241 -1597 2341 -1581
rect 2399 -1547 2499 -1500
rect 2399 -1581 2415 -1547
rect 2483 -1581 2499 -1547
rect 2399 -1597 2499 -1581
rect 2557 -1547 2657 -1500
rect 2557 -1581 2573 -1547
rect 2641 -1581 2657 -1547
rect 2557 -1597 2657 -1581
rect 2715 -1547 2815 -1500
rect 2715 -1581 2731 -1547
rect 2799 -1581 2815 -1547
rect 2715 -1597 2815 -1581
rect 2873 -1547 2973 -1500
rect 2873 -1581 2889 -1547
rect 2957 -1581 2973 -1547
rect 2873 -1597 2973 -1581
rect 3031 -1547 3131 -1500
rect 3031 -1581 3047 -1547
rect 3115 -1581 3131 -1547
rect 3031 -1597 3131 -1581
rect 3189 -1547 3289 -1500
rect 3189 -1581 3205 -1547
rect 3273 -1581 3289 -1547
rect 3189 -1597 3289 -1581
rect 3347 -1547 3447 -1500
rect 3347 -1581 3363 -1547
rect 3431 -1581 3447 -1547
rect 3347 -1597 3447 -1581
rect 3505 -1547 3605 -1500
rect 3505 -1581 3521 -1547
rect 3589 -1581 3605 -1547
rect 3505 -1597 3605 -1581
rect 3663 -1547 3763 -1500
rect 3663 -1581 3679 -1547
rect 3747 -1581 3763 -1547
rect 3663 -1597 3763 -1581
rect 3821 -1547 3921 -1500
rect 3821 -1581 3837 -1547
rect 3905 -1581 3921 -1547
rect 3821 -1597 3921 -1581
rect 3979 -1547 4079 -1500
rect 3979 -1581 3995 -1547
rect 4063 -1581 4079 -1547
rect 3979 -1597 4079 -1581
rect 4137 -1547 4237 -1500
rect 4137 -1581 4153 -1547
rect 4221 -1581 4237 -1547
rect 4137 -1597 4237 -1581
rect 4295 -1547 4395 -1500
rect 4295 -1581 4311 -1547
rect 4379 -1581 4395 -1547
rect 4295 -1597 4395 -1581
rect 4453 -1547 4553 -1500
rect 4453 -1581 4469 -1547
rect 4537 -1581 4553 -1547
rect 4453 -1597 4553 -1581
rect 4611 -1547 4711 -1500
rect 4611 -1581 4627 -1547
rect 4695 -1581 4711 -1547
rect 4611 -1597 4711 -1581
rect 4769 -1547 4869 -1500
rect 4769 -1581 4785 -1547
rect 4853 -1581 4869 -1547
rect 4769 -1597 4869 -1581
rect 4927 -1547 5027 -1500
rect 4927 -1581 4943 -1547
rect 5011 -1581 5027 -1547
rect 4927 -1597 5027 -1581
rect 5085 -1547 5185 -1500
rect 5085 -1581 5101 -1547
rect 5169 -1581 5185 -1547
rect 5085 -1597 5185 -1581
rect 5243 -1547 5343 -1500
rect 5243 -1581 5259 -1547
rect 5327 -1581 5343 -1547
rect 5243 -1597 5343 -1581
rect 5401 -1547 5501 -1500
rect 5401 -1581 5417 -1547
rect 5485 -1581 5501 -1547
rect 5401 -1597 5501 -1581
rect 5559 -1547 5659 -1500
rect 5559 -1581 5575 -1547
rect 5643 -1581 5659 -1547
rect 5559 -1597 5659 -1581
rect 5717 -1547 5817 -1500
rect 5717 -1581 5733 -1547
rect 5801 -1581 5817 -1547
rect 5717 -1597 5817 -1581
rect 5875 -1547 5975 -1500
rect 5875 -1581 5891 -1547
rect 5959 -1581 5975 -1547
rect 5875 -1597 5975 -1581
rect 6033 -1547 6133 -1500
rect 6033 -1581 6049 -1547
rect 6117 -1581 6133 -1547
rect 6033 -1597 6133 -1581
rect 6191 -1547 6291 -1500
rect 6191 -1581 6207 -1547
rect 6275 -1581 6291 -1547
rect 6191 -1597 6291 -1581
rect 6349 -1547 6449 -1500
rect 6349 -1581 6365 -1547
rect 6433 -1581 6449 -1547
rect 6349 -1597 6449 -1581
rect 6507 -1547 6607 -1500
rect 6507 -1581 6523 -1547
rect 6591 -1581 6607 -1547
rect 6507 -1597 6607 -1581
rect 6665 -1547 6765 -1500
rect 6665 -1581 6681 -1547
rect 6749 -1581 6765 -1547
rect 6665 -1597 6765 -1581
rect 6823 -1547 6923 -1500
rect 6823 -1581 6839 -1547
rect 6907 -1581 6923 -1547
rect 6823 -1597 6923 -1581
<< polycont >>
rect -6907 1547 -6839 1581
rect -6749 1547 -6681 1581
rect -6591 1547 -6523 1581
rect -6433 1547 -6365 1581
rect -6275 1547 -6207 1581
rect -6117 1547 -6049 1581
rect -5959 1547 -5891 1581
rect -5801 1547 -5733 1581
rect -5643 1547 -5575 1581
rect -5485 1547 -5417 1581
rect -5327 1547 -5259 1581
rect -5169 1547 -5101 1581
rect -5011 1547 -4943 1581
rect -4853 1547 -4785 1581
rect -4695 1547 -4627 1581
rect -4537 1547 -4469 1581
rect -4379 1547 -4311 1581
rect -4221 1547 -4153 1581
rect -4063 1547 -3995 1581
rect -3905 1547 -3837 1581
rect -3747 1547 -3679 1581
rect -3589 1547 -3521 1581
rect -3431 1547 -3363 1581
rect -3273 1547 -3205 1581
rect -3115 1547 -3047 1581
rect -2957 1547 -2889 1581
rect -2799 1547 -2731 1581
rect -2641 1547 -2573 1581
rect -2483 1547 -2415 1581
rect -2325 1547 -2257 1581
rect -2167 1547 -2099 1581
rect -2009 1547 -1941 1581
rect -1851 1547 -1783 1581
rect -1693 1547 -1625 1581
rect -1535 1547 -1467 1581
rect -1377 1547 -1309 1581
rect -1219 1547 -1151 1581
rect -1061 1547 -993 1581
rect -903 1547 -835 1581
rect -745 1547 -677 1581
rect -587 1547 -519 1581
rect -429 1547 -361 1581
rect -271 1547 -203 1581
rect -113 1547 -45 1581
rect 45 1547 113 1581
rect 203 1547 271 1581
rect 361 1547 429 1581
rect 519 1547 587 1581
rect 677 1547 745 1581
rect 835 1547 903 1581
rect 993 1547 1061 1581
rect 1151 1547 1219 1581
rect 1309 1547 1377 1581
rect 1467 1547 1535 1581
rect 1625 1547 1693 1581
rect 1783 1547 1851 1581
rect 1941 1547 2009 1581
rect 2099 1547 2167 1581
rect 2257 1547 2325 1581
rect 2415 1547 2483 1581
rect 2573 1547 2641 1581
rect 2731 1547 2799 1581
rect 2889 1547 2957 1581
rect 3047 1547 3115 1581
rect 3205 1547 3273 1581
rect 3363 1547 3431 1581
rect 3521 1547 3589 1581
rect 3679 1547 3747 1581
rect 3837 1547 3905 1581
rect 3995 1547 4063 1581
rect 4153 1547 4221 1581
rect 4311 1547 4379 1581
rect 4469 1547 4537 1581
rect 4627 1547 4695 1581
rect 4785 1547 4853 1581
rect 4943 1547 5011 1581
rect 5101 1547 5169 1581
rect 5259 1547 5327 1581
rect 5417 1547 5485 1581
rect 5575 1547 5643 1581
rect 5733 1547 5801 1581
rect 5891 1547 5959 1581
rect 6049 1547 6117 1581
rect 6207 1547 6275 1581
rect 6365 1547 6433 1581
rect 6523 1547 6591 1581
rect 6681 1547 6749 1581
rect 6839 1547 6907 1581
rect -6907 -1581 -6839 -1547
rect -6749 -1581 -6681 -1547
rect -6591 -1581 -6523 -1547
rect -6433 -1581 -6365 -1547
rect -6275 -1581 -6207 -1547
rect -6117 -1581 -6049 -1547
rect -5959 -1581 -5891 -1547
rect -5801 -1581 -5733 -1547
rect -5643 -1581 -5575 -1547
rect -5485 -1581 -5417 -1547
rect -5327 -1581 -5259 -1547
rect -5169 -1581 -5101 -1547
rect -5011 -1581 -4943 -1547
rect -4853 -1581 -4785 -1547
rect -4695 -1581 -4627 -1547
rect -4537 -1581 -4469 -1547
rect -4379 -1581 -4311 -1547
rect -4221 -1581 -4153 -1547
rect -4063 -1581 -3995 -1547
rect -3905 -1581 -3837 -1547
rect -3747 -1581 -3679 -1547
rect -3589 -1581 -3521 -1547
rect -3431 -1581 -3363 -1547
rect -3273 -1581 -3205 -1547
rect -3115 -1581 -3047 -1547
rect -2957 -1581 -2889 -1547
rect -2799 -1581 -2731 -1547
rect -2641 -1581 -2573 -1547
rect -2483 -1581 -2415 -1547
rect -2325 -1581 -2257 -1547
rect -2167 -1581 -2099 -1547
rect -2009 -1581 -1941 -1547
rect -1851 -1581 -1783 -1547
rect -1693 -1581 -1625 -1547
rect -1535 -1581 -1467 -1547
rect -1377 -1581 -1309 -1547
rect -1219 -1581 -1151 -1547
rect -1061 -1581 -993 -1547
rect -903 -1581 -835 -1547
rect -745 -1581 -677 -1547
rect -587 -1581 -519 -1547
rect -429 -1581 -361 -1547
rect -271 -1581 -203 -1547
rect -113 -1581 -45 -1547
rect 45 -1581 113 -1547
rect 203 -1581 271 -1547
rect 361 -1581 429 -1547
rect 519 -1581 587 -1547
rect 677 -1581 745 -1547
rect 835 -1581 903 -1547
rect 993 -1581 1061 -1547
rect 1151 -1581 1219 -1547
rect 1309 -1581 1377 -1547
rect 1467 -1581 1535 -1547
rect 1625 -1581 1693 -1547
rect 1783 -1581 1851 -1547
rect 1941 -1581 2009 -1547
rect 2099 -1581 2167 -1547
rect 2257 -1581 2325 -1547
rect 2415 -1581 2483 -1547
rect 2573 -1581 2641 -1547
rect 2731 -1581 2799 -1547
rect 2889 -1581 2957 -1547
rect 3047 -1581 3115 -1547
rect 3205 -1581 3273 -1547
rect 3363 -1581 3431 -1547
rect 3521 -1581 3589 -1547
rect 3679 -1581 3747 -1547
rect 3837 -1581 3905 -1547
rect 3995 -1581 4063 -1547
rect 4153 -1581 4221 -1547
rect 4311 -1581 4379 -1547
rect 4469 -1581 4537 -1547
rect 4627 -1581 4695 -1547
rect 4785 -1581 4853 -1547
rect 4943 -1581 5011 -1547
rect 5101 -1581 5169 -1547
rect 5259 -1581 5327 -1547
rect 5417 -1581 5485 -1547
rect 5575 -1581 5643 -1547
rect 5733 -1581 5801 -1547
rect 5891 -1581 5959 -1547
rect 6049 -1581 6117 -1547
rect 6207 -1581 6275 -1547
rect 6365 -1581 6433 -1547
rect 6523 -1581 6591 -1547
rect 6681 -1581 6749 -1547
rect 6839 -1581 6907 -1547
<< locali >>
rect -6923 1547 -6907 1581
rect -6839 1547 -6823 1581
rect -6765 1547 -6749 1581
rect -6681 1547 -6665 1581
rect -6607 1547 -6591 1581
rect -6523 1547 -6507 1581
rect -6449 1547 -6433 1581
rect -6365 1547 -6349 1581
rect -6291 1547 -6275 1581
rect -6207 1547 -6191 1581
rect -6133 1547 -6117 1581
rect -6049 1547 -6033 1581
rect -5975 1547 -5959 1581
rect -5891 1547 -5875 1581
rect -5817 1547 -5801 1581
rect -5733 1547 -5717 1581
rect -5659 1547 -5643 1581
rect -5575 1547 -5559 1581
rect -5501 1547 -5485 1581
rect -5417 1547 -5401 1581
rect -5343 1547 -5327 1581
rect -5259 1547 -5243 1581
rect -5185 1547 -5169 1581
rect -5101 1547 -5085 1581
rect -5027 1547 -5011 1581
rect -4943 1547 -4927 1581
rect -4869 1547 -4853 1581
rect -4785 1547 -4769 1581
rect -4711 1547 -4695 1581
rect -4627 1547 -4611 1581
rect -4553 1547 -4537 1581
rect -4469 1547 -4453 1581
rect -4395 1547 -4379 1581
rect -4311 1547 -4295 1581
rect -4237 1547 -4221 1581
rect -4153 1547 -4137 1581
rect -4079 1547 -4063 1581
rect -3995 1547 -3979 1581
rect -3921 1547 -3905 1581
rect -3837 1547 -3821 1581
rect -3763 1547 -3747 1581
rect -3679 1547 -3663 1581
rect -3605 1547 -3589 1581
rect -3521 1547 -3505 1581
rect -3447 1547 -3431 1581
rect -3363 1547 -3347 1581
rect -3289 1547 -3273 1581
rect -3205 1547 -3189 1581
rect -3131 1547 -3115 1581
rect -3047 1547 -3031 1581
rect -2973 1547 -2957 1581
rect -2889 1547 -2873 1581
rect -2815 1547 -2799 1581
rect -2731 1547 -2715 1581
rect -2657 1547 -2641 1581
rect -2573 1547 -2557 1581
rect -2499 1547 -2483 1581
rect -2415 1547 -2399 1581
rect -2341 1547 -2325 1581
rect -2257 1547 -2241 1581
rect -2183 1547 -2167 1581
rect -2099 1547 -2083 1581
rect -2025 1547 -2009 1581
rect -1941 1547 -1925 1581
rect -1867 1547 -1851 1581
rect -1783 1547 -1767 1581
rect -1709 1547 -1693 1581
rect -1625 1547 -1609 1581
rect -1551 1547 -1535 1581
rect -1467 1547 -1451 1581
rect -1393 1547 -1377 1581
rect -1309 1547 -1293 1581
rect -1235 1547 -1219 1581
rect -1151 1547 -1135 1581
rect -1077 1547 -1061 1581
rect -993 1547 -977 1581
rect -919 1547 -903 1581
rect -835 1547 -819 1581
rect -761 1547 -745 1581
rect -677 1547 -661 1581
rect -603 1547 -587 1581
rect -519 1547 -503 1581
rect -445 1547 -429 1581
rect -361 1547 -345 1581
rect -287 1547 -271 1581
rect -203 1547 -187 1581
rect -129 1547 -113 1581
rect -45 1547 -29 1581
rect 29 1547 45 1581
rect 113 1547 129 1581
rect 187 1547 203 1581
rect 271 1547 287 1581
rect 345 1547 361 1581
rect 429 1547 445 1581
rect 503 1547 519 1581
rect 587 1547 603 1581
rect 661 1547 677 1581
rect 745 1547 761 1581
rect 819 1547 835 1581
rect 903 1547 919 1581
rect 977 1547 993 1581
rect 1061 1547 1077 1581
rect 1135 1547 1151 1581
rect 1219 1547 1235 1581
rect 1293 1547 1309 1581
rect 1377 1547 1393 1581
rect 1451 1547 1467 1581
rect 1535 1547 1551 1581
rect 1609 1547 1625 1581
rect 1693 1547 1709 1581
rect 1767 1547 1783 1581
rect 1851 1547 1867 1581
rect 1925 1547 1941 1581
rect 2009 1547 2025 1581
rect 2083 1547 2099 1581
rect 2167 1547 2183 1581
rect 2241 1547 2257 1581
rect 2325 1547 2341 1581
rect 2399 1547 2415 1581
rect 2483 1547 2499 1581
rect 2557 1547 2573 1581
rect 2641 1547 2657 1581
rect 2715 1547 2731 1581
rect 2799 1547 2815 1581
rect 2873 1547 2889 1581
rect 2957 1547 2973 1581
rect 3031 1547 3047 1581
rect 3115 1547 3131 1581
rect 3189 1547 3205 1581
rect 3273 1547 3289 1581
rect 3347 1547 3363 1581
rect 3431 1547 3447 1581
rect 3505 1547 3521 1581
rect 3589 1547 3605 1581
rect 3663 1547 3679 1581
rect 3747 1547 3763 1581
rect 3821 1547 3837 1581
rect 3905 1547 3921 1581
rect 3979 1547 3995 1581
rect 4063 1547 4079 1581
rect 4137 1547 4153 1581
rect 4221 1547 4237 1581
rect 4295 1547 4311 1581
rect 4379 1547 4395 1581
rect 4453 1547 4469 1581
rect 4537 1547 4553 1581
rect 4611 1547 4627 1581
rect 4695 1547 4711 1581
rect 4769 1547 4785 1581
rect 4853 1547 4869 1581
rect 4927 1547 4943 1581
rect 5011 1547 5027 1581
rect 5085 1547 5101 1581
rect 5169 1547 5185 1581
rect 5243 1547 5259 1581
rect 5327 1547 5343 1581
rect 5401 1547 5417 1581
rect 5485 1547 5501 1581
rect 5559 1547 5575 1581
rect 5643 1547 5659 1581
rect 5717 1547 5733 1581
rect 5801 1547 5817 1581
rect 5875 1547 5891 1581
rect 5959 1547 5975 1581
rect 6033 1547 6049 1581
rect 6117 1547 6133 1581
rect 6191 1547 6207 1581
rect 6275 1547 6291 1581
rect 6349 1547 6365 1581
rect 6433 1547 6449 1581
rect 6507 1547 6523 1581
rect 6591 1547 6607 1581
rect 6665 1547 6681 1581
rect 6749 1547 6765 1581
rect 6823 1547 6839 1581
rect 6907 1547 6923 1581
rect -6969 1488 -6935 1504
rect -6969 -1504 -6935 -1488
rect -6811 1488 -6777 1504
rect -6811 -1504 -6777 -1488
rect -6653 1488 -6619 1504
rect -6653 -1504 -6619 -1488
rect -6495 1488 -6461 1504
rect -6495 -1504 -6461 -1488
rect -6337 1488 -6303 1504
rect -6337 -1504 -6303 -1488
rect -6179 1488 -6145 1504
rect -6179 -1504 -6145 -1488
rect -6021 1488 -5987 1504
rect -6021 -1504 -5987 -1488
rect -5863 1488 -5829 1504
rect -5863 -1504 -5829 -1488
rect -5705 1488 -5671 1504
rect -5705 -1504 -5671 -1488
rect -5547 1488 -5513 1504
rect -5547 -1504 -5513 -1488
rect -5389 1488 -5355 1504
rect -5389 -1504 -5355 -1488
rect -5231 1488 -5197 1504
rect -5231 -1504 -5197 -1488
rect -5073 1488 -5039 1504
rect -5073 -1504 -5039 -1488
rect -4915 1488 -4881 1504
rect -4915 -1504 -4881 -1488
rect -4757 1488 -4723 1504
rect -4757 -1504 -4723 -1488
rect -4599 1488 -4565 1504
rect -4599 -1504 -4565 -1488
rect -4441 1488 -4407 1504
rect -4441 -1504 -4407 -1488
rect -4283 1488 -4249 1504
rect -4283 -1504 -4249 -1488
rect -4125 1488 -4091 1504
rect -4125 -1504 -4091 -1488
rect -3967 1488 -3933 1504
rect -3967 -1504 -3933 -1488
rect -3809 1488 -3775 1504
rect -3809 -1504 -3775 -1488
rect -3651 1488 -3617 1504
rect -3651 -1504 -3617 -1488
rect -3493 1488 -3459 1504
rect -3493 -1504 -3459 -1488
rect -3335 1488 -3301 1504
rect -3335 -1504 -3301 -1488
rect -3177 1488 -3143 1504
rect -3177 -1504 -3143 -1488
rect -3019 1488 -2985 1504
rect -3019 -1504 -2985 -1488
rect -2861 1488 -2827 1504
rect -2861 -1504 -2827 -1488
rect -2703 1488 -2669 1504
rect -2703 -1504 -2669 -1488
rect -2545 1488 -2511 1504
rect -2545 -1504 -2511 -1488
rect -2387 1488 -2353 1504
rect -2387 -1504 -2353 -1488
rect -2229 1488 -2195 1504
rect -2229 -1504 -2195 -1488
rect -2071 1488 -2037 1504
rect -2071 -1504 -2037 -1488
rect -1913 1488 -1879 1504
rect -1913 -1504 -1879 -1488
rect -1755 1488 -1721 1504
rect -1755 -1504 -1721 -1488
rect -1597 1488 -1563 1504
rect -1597 -1504 -1563 -1488
rect -1439 1488 -1405 1504
rect -1439 -1504 -1405 -1488
rect -1281 1488 -1247 1504
rect -1281 -1504 -1247 -1488
rect -1123 1488 -1089 1504
rect -1123 -1504 -1089 -1488
rect -965 1488 -931 1504
rect -965 -1504 -931 -1488
rect -807 1488 -773 1504
rect -807 -1504 -773 -1488
rect -649 1488 -615 1504
rect -649 -1504 -615 -1488
rect -491 1488 -457 1504
rect -491 -1504 -457 -1488
rect -333 1488 -299 1504
rect -333 -1504 -299 -1488
rect -175 1488 -141 1504
rect -175 -1504 -141 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 141 1488 175 1504
rect 141 -1504 175 -1488
rect 299 1488 333 1504
rect 299 -1504 333 -1488
rect 457 1488 491 1504
rect 457 -1504 491 -1488
rect 615 1488 649 1504
rect 615 -1504 649 -1488
rect 773 1488 807 1504
rect 773 -1504 807 -1488
rect 931 1488 965 1504
rect 931 -1504 965 -1488
rect 1089 1488 1123 1504
rect 1089 -1504 1123 -1488
rect 1247 1488 1281 1504
rect 1247 -1504 1281 -1488
rect 1405 1488 1439 1504
rect 1405 -1504 1439 -1488
rect 1563 1488 1597 1504
rect 1563 -1504 1597 -1488
rect 1721 1488 1755 1504
rect 1721 -1504 1755 -1488
rect 1879 1488 1913 1504
rect 1879 -1504 1913 -1488
rect 2037 1488 2071 1504
rect 2037 -1504 2071 -1488
rect 2195 1488 2229 1504
rect 2195 -1504 2229 -1488
rect 2353 1488 2387 1504
rect 2353 -1504 2387 -1488
rect 2511 1488 2545 1504
rect 2511 -1504 2545 -1488
rect 2669 1488 2703 1504
rect 2669 -1504 2703 -1488
rect 2827 1488 2861 1504
rect 2827 -1504 2861 -1488
rect 2985 1488 3019 1504
rect 2985 -1504 3019 -1488
rect 3143 1488 3177 1504
rect 3143 -1504 3177 -1488
rect 3301 1488 3335 1504
rect 3301 -1504 3335 -1488
rect 3459 1488 3493 1504
rect 3459 -1504 3493 -1488
rect 3617 1488 3651 1504
rect 3617 -1504 3651 -1488
rect 3775 1488 3809 1504
rect 3775 -1504 3809 -1488
rect 3933 1488 3967 1504
rect 3933 -1504 3967 -1488
rect 4091 1488 4125 1504
rect 4091 -1504 4125 -1488
rect 4249 1488 4283 1504
rect 4249 -1504 4283 -1488
rect 4407 1488 4441 1504
rect 4407 -1504 4441 -1488
rect 4565 1488 4599 1504
rect 4565 -1504 4599 -1488
rect 4723 1488 4757 1504
rect 4723 -1504 4757 -1488
rect 4881 1488 4915 1504
rect 4881 -1504 4915 -1488
rect 5039 1488 5073 1504
rect 5039 -1504 5073 -1488
rect 5197 1488 5231 1504
rect 5197 -1504 5231 -1488
rect 5355 1488 5389 1504
rect 5355 -1504 5389 -1488
rect 5513 1488 5547 1504
rect 5513 -1504 5547 -1488
rect 5671 1488 5705 1504
rect 5671 -1504 5705 -1488
rect 5829 1488 5863 1504
rect 5829 -1504 5863 -1488
rect 5987 1488 6021 1504
rect 5987 -1504 6021 -1488
rect 6145 1488 6179 1504
rect 6145 -1504 6179 -1488
rect 6303 1488 6337 1504
rect 6303 -1504 6337 -1488
rect 6461 1488 6495 1504
rect 6461 -1504 6495 -1488
rect 6619 1488 6653 1504
rect 6619 -1504 6653 -1488
rect 6777 1488 6811 1504
rect 6777 -1504 6811 -1488
rect 6935 1488 6969 1504
rect 6935 -1504 6969 -1488
rect -6923 -1581 -6907 -1547
rect -6839 -1581 -6823 -1547
rect -6765 -1581 -6749 -1547
rect -6681 -1581 -6665 -1547
rect -6607 -1581 -6591 -1547
rect -6523 -1581 -6507 -1547
rect -6449 -1581 -6433 -1547
rect -6365 -1581 -6349 -1547
rect -6291 -1581 -6275 -1547
rect -6207 -1581 -6191 -1547
rect -6133 -1581 -6117 -1547
rect -6049 -1581 -6033 -1547
rect -5975 -1581 -5959 -1547
rect -5891 -1581 -5875 -1547
rect -5817 -1581 -5801 -1547
rect -5733 -1581 -5717 -1547
rect -5659 -1581 -5643 -1547
rect -5575 -1581 -5559 -1547
rect -5501 -1581 -5485 -1547
rect -5417 -1581 -5401 -1547
rect -5343 -1581 -5327 -1547
rect -5259 -1581 -5243 -1547
rect -5185 -1581 -5169 -1547
rect -5101 -1581 -5085 -1547
rect -5027 -1581 -5011 -1547
rect -4943 -1581 -4927 -1547
rect -4869 -1581 -4853 -1547
rect -4785 -1581 -4769 -1547
rect -4711 -1581 -4695 -1547
rect -4627 -1581 -4611 -1547
rect -4553 -1581 -4537 -1547
rect -4469 -1581 -4453 -1547
rect -4395 -1581 -4379 -1547
rect -4311 -1581 -4295 -1547
rect -4237 -1581 -4221 -1547
rect -4153 -1581 -4137 -1547
rect -4079 -1581 -4063 -1547
rect -3995 -1581 -3979 -1547
rect -3921 -1581 -3905 -1547
rect -3837 -1581 -3821 -1547
rect -3763 -1581 -3747 -1547
rect -3679 -1581 -3663 -1547
rect -3605 -1581 -3589 -1547
rect -3521 -1581 -3505 -1547
rect -3447 -1581 -3431 -1547
rect -3363 -1581 -3347 -1547
rect -3289 -1581 -3273 -1547
rect -3205 -1581 -3189 -1547
rect -3131 -1581 -3115 -1547
rect -3047 -1581 -3031 -1547
rect -2973 -1581 -2957 -1547
rect -2889 -1581 -2873 -1547
rect -2815 -1581 -2799 -1547
rect -2731 -1581 -2715 -1547
rect -2657 -1581 -2641 -1547
rect -2573 -1581 -2557 -1547
rect -2499 -1581 -2483 -1547
rect -2415 -1581 -2399 -1547
rect -2341 -1581 -2325 -1547
rect -2257 -1581 -2241 -1547
rect -2183 -1581 -2167 -1547
rect -2099 -1581 -2083 -1547
rect -2025 -1581 -2009 -1547
rect -1941 -1581 -1925 -1547
rect -1867 -1581 -1851 -1547
rect -1783 -1581 -1767 -1547
rect -1709 -1581 -1693 -1547
rect -1625 -1581 -1609 -1547
rect -1551 -1581 -1535 -1547
rect -1467 -1581 -1451 -1547
rect -1393 -1581 -1377 -1547
rect -1309 -1581 -1293 -1547
rect -1235 -1581 -1219 -1547
rect -1151 -1581 -1135 -1547
rect -1077 -1581 -1061 -1547
rect -993 -1581 -977 -1547
rect -919 -1581 -903 -1547
rect -835 -1581 -819 -1547
rect -761 -1581 -745 -1547
rect -677 -1581 -661 -1547
rect -603 -1581 -587 -1547
rect -519 -1581 -503 -1547
rect -445 -1581 -429 -1547
rect -361 -1581 -345 -1547
rect -287 -1581 -271 -1547
rect -203 -1581 -187 -1547
rect -129 -1581 -113 -1547
rect -45 -1581 -29 -1547
rect 29 -1581 45 -1547
rect 113 -1581 129 -1547
rect 187 -1581 203 -1547
rect 271 -1581 287 -1547
rect 345 -1581 361 -1547
rect 429 -1581 445 -1547
rect 503 -1581 519 -1547
rect 587 -1581 603 -1547
rect 661 -1581 677 -1547
rect 745 -1581 761 -1547
rect 819 -1581 835 -1547
rect 903 -1581 919 -1547
rect 977 -1581 993 -1547
rect 1061 -1581 1077 -1547
rect 1135 -1581 1151 -1547
rect 1219 -1581 1235 -1547
rect 1293 -1581 1309 -1547
rect 1377 -1581 1393 -1547
rect 1451 -1581 1467 -1547
rect 1535 -1581 1551 -1547
rect 1609 -1581 1625 -1547
rect 1693 -1581 1709 -1547
rect 1767 -1581 1783 -1547
rect 1851 -1581 1867 -1547
rect 1925 -1581 1941 -1547
rect 2009 -1581 2025 -1547
rect 2083 -1581 2099 -1547
rect 2167 -1581 2183 -1547
rect 2241 -1581 2257 -1547
rect 2325 -1581 2341 -1547
rect 2399 -1581 2415 -1547
rect 2483 -1581 2499 -1547
rect 2557 -1581 2573 -1547
rect 2641 -1581 2657 -1547
rect 2715 -1581 2731 -1547
rect 2799 -1581 2815 -1547
rect 2873 -1581 2889 -1547
rect 2957 -1581 2973 -1547
rect 3031 -1581 3047 -1547
rect 3115 -1581 3131 -1547
rect 3189 -1581 3205 -1547
rect 3273 -1581 3289 -1547
rect 3347 -1581 3363 -1547
rect 3431 -1581 3447 -1547
rect 3505 -1581 3521 -1547
rect 3589 -1581 3605 -1547
rect 3663 -1581 3679 -1547
rect 3747 -1581 3763 -1547
rect 3821 -1581 3837 -1547
rect 3905 -1581 3921 -1547
rect 3979 -1581 3995 -1547
rect 4063 -1581 4079 -1547
rect 4137 -1581 4153 -1547
rect 4221 -1581 4237 -1547
rect 4295 -1581 4311 -1547
rect 4379 -1581 4395 -1547
rect 4453 -1581 4469 -1547
rect 4537 -1581 4553 -1547
rect 4611 -1581 4627 -1547
rect 4695 -1581 4711 -1547
rect 4769 -1581 4785 -1547
rect 4853 -1581 4869 -1547
rect 4927 -1581 4943 -1547
rect 5011 -1581 5027 -1547
rect 5085 -1581 5101 -1547
rect 5169 -1581 5185 -1547
rect 5243 -1581 5259 -1547
rect 5327 -1581 5343 -1547
rect 5401 -1581 5417 -1547
rect 5485 -1581 5501 -1547
rect 5559 -1581 5575 -1547
rect 5643 -1581 5659 -1547
rect 5717 -1581 5733 -1547
rect 5801 -1581 5817 -1547
rect 5875 -1581 5891 -1547
rect 5959 -1581 5975 -1547
rect 6033 -1581 6049 -1547
rect 6117 -1581 6133 -1547
rect 6191 -1581 6207 -1547
rect 6275 -1581 6291 -1547
rect 6349 -1581 6365 -1547
rect 6433 -1581 6449 -1547
rect 6507 -1581 6523 -1547
rect 6591 -1581 6607 -1547
rect 6665 -1581 6681 -1547
rect 6749 -1581 6765 -1547
rect 6823 -1581 6839 -1547
rect 6907 -1581 6923 -1547
<< viali >>
rect -6969 -1488 -6935 1488
rect -6811 -1488 -6777 1488
rect -6653 -1488 -6619 1488
rect -6495 -1488 -6461 1488
rect -6337 -1488 -6303 1488
rect -6179 -1488 -6145 1488
rect -6021 -1488 -5987 1488
rect -5863 -1488 -5829 1488
rect -5705 -1488 -5671 1488
rect -5547 -1488 -5513 1488
rect -5389 -1488 -5355 1488
rect -5231 -1488 -5197 1488
rect -5073 -1488 -5039 1488
rect -4915 -1488 -4881 1488
rect -4757 -1488 -4723 1488
rect -4599 -1488 -4565 1488
rect -4441 -1488 -4407 1488
rect -4283 -1488 -4249 1488
rect -4125 -1488 -4091 1488
rect -3967 -1488 -3933 1488
rect -3809 -1488 -3775 1488
rect -3651 -1488 -3617 1488
rect -3493 -1488 -3459 1488
rect -3335 -1488 -3301 1488
rect -3177 -1488 -3143 1488
rect -3019 -1488 -2985 1488
rect -2861 -1488 -2827 1488
rect -2703 -1488 -2669 1488
rect -2545 -1488 -2511 1488
rect -2387 -1488 -2353 1488
rect -2229 -1488 -2195 1488
rect -2071 -1488 -2037 1488
rect -1913 -1488 -1879 1488
rect -1755 -1488 -1721 1488
rect -1597 -1488 -1563 1488
rect -1439 -1488 -1405 1488
rect -1281 -1488 -1247 1488
rect -1123 -1488 -1089 1488
rect -965 -1488 -931 1488
rect -807 -1488 -773 1488
rect -649 -1488 -615 1488
rect -491 -1488 -457 1488
rect -333 -1488 -299 1488
rect -175 -1488 -141 1488
rect -17 -1488 17 1488
rect 141 -1488 175 1488
rect 299 -1488 333 1488
rect 457 -1488 491 1488
rect 615 -1488 649 1488
rect 773 -1488 807 1488
rect 931 -1488 965 1488
rect 1089 -1488 1123 1488
rect 1247 -1488 1281 1488
rect 1405 -1488 1439 1488
rect 1563 -1488 1597 1488
rect 1721 -1488 1755 1488
rect 1879 -1488 1913 1488
rect 2037 -1488 2071 1488
rect 2195 -1488 2229 1488
rect 2353 -1488 2387 1488
rect 2511 -1488 2545 1488
rect 2669 -1488 2703 1488
rect 2827 -1488 2861 1488
rect 2985 -1488 3019 1488
rect 3143 -1488 3177 1488
rect 3301 -1488 3335 1488
rect 3459 -1488 3493 1488
rect 3617 -1488 3651 1488
rect 3775 -1488 3809 1488
rect 3933 -1488 3967 1488
rect 4091 -1488 4125 1488
rect 4249 -1488 4283 1488
rect 4407 -1488 4441 1488
rect 4565 -1488 4599 1488
rect 4723 -1488 4757 1488
rect 4881 -1488 4915 1488
rect 5039 -1488 5073 1488
rect 5197 -1488 5231 1488
rect 5355 -1488 5389 1488
rect 5513 -1488 5547 1488
rect 5671 -1488 5705 1488
rect 5829 -1488 5863 1488
rect 5987 -1488 6021 1488
rect 6145 -1488 6179 1488
rect 6303 -1488 6337 1488
rect 6461 -1488 6495 1488
rect 6619 -1488 6653 1488
rect 6777 -1488 6811 1488
rect 6935 -1488 6969 1488
<< metal1 >>
rect -6975 1488 -6929 1500
rect -6975 -1488 -6969 1488
rect -6935 -1488 -6929 1488
rect -6975 -1500 -6929 -1488
rect -6817 1488 -6771 1500
rect -6817 -1488 -6811 1488
rect -6777 -1488 -6771 1488
rect -6817 -1500 -6771 -1488
rect -6659 1488 -6613 1500
rect -6659 -1488 -6653 1488
rect -6619 -1488 -6613 1488
rect -6659 -1500 -6613 -1488
rect -6501 1488 -6455 1500
rect -6501 -1488 -6495 1488
rect -6461 -1488 -6455 1488
rect -6501 -1500 -6455 -1488
rect -6343 1488 -6297 1500
rect -6343 -1488 -6337 1488
rect -6303 -1488 -6297 1488
rect -6343 -1500 -6297 -1488
rect -6185 1488 -6139 1500
rect -6185 -1488 -6179 1488
rect -6145 -1488 -6139 1488
rect -6185 -1500 -6139 -1488
rect -6027 1488 -5981 1500
rect -6027 -1488 -6021 1488
rect -5987 -1488 -5981 1488
rect -6027 -1500 -5981 -1488
rect -5869 1488 -5823 1500
rect -5869 -1488 -5863 1488
rect -5829 -1488 -5823 1488
rect -5869 -1500 -5823 -1488
rect -5711 1488 -5665 1500
rect -5711 -1488 -5705 1488
rect -5671 -1488 -5665 1488
rect -5711 -1500 -5665 -1488
rect -5553 1488 -5507 1500
rect -5553 -1488 -5547 1488
rect -5513 -1488 -5507 1488
rect -5553 -1500 -5507 -1488
rect -5395 1488 -5349 1500
rect -5395 -1488 -5389 1488
rect -5355 -1488 -5349 1488
rect -5395 -1500 -5349 -1488
rect -5237 1488 -5191 1500
rect -5237 -1488 -5231 1488
rect -5197 -1488 -5191 1488
rect -5237 -1500 -5191 -1488
rect -5079 1488 -5033 1500
rect -5079 -1488 -5073 1488
rect -5039 -1488 -5033 1488
rect -5079 -1500 -5033 -1488
rect -4921 1488 -4875 1500
rect -4921 -1488 -4915 1488
rect -4881 -1488 -4875 1488
rect -4921 -1500 -4875 -1488
rect -4763 1488 -4717 1500
rect -4763 -1488 -4757 1488
rect -4723 -1488 -4717 1488
rect -4763 -1500 -4717 -1488
rect -4605 1488 -4559 1500
rect -4605 -1488 -4599 1488
rect -4565 -1488 -4559 1488
rect -4605 -1500 -4559 -1488
rect -4447 1488 -4401 1500
rect -4447 -1488 -4441 1488
rect -4407 -1488 -4401 1488
rect -4447 -1500 -4401 -1488
rect -4289 1488 -4243 1500
rect -4289 -1488 -4283 1488
rect -4249 -1488 -4243 1488
rect -4289 -1500 -4243 -1488
rect -4131 1488 -4085 1500
rect -4131 -1488 -4125 1488
rect -4091 -1488 -4085 1488
rect -4131 -1500 -4085 -1488
rect -3973 1488 -3927 1500
rect -3973 -1488 -3967 1488
rect -3933 -1488 -3927 1488
rect -3973 -1500 -3927 -1488
rect -3815 1488 -3769 1500
rect -3815 -1488 -3809 1488
rect -3775 -1488 -3769 1488
rect -3815 -1500 -3769 -1488
rect -3657 1488 -3611 1500
rect -3657 -1488 -3651 1488
rect -3617 -1488 -3611 1488
rect -3657 -1500 -3611 -1488
rect -3499 1488 -3453 1500
rect -3499 -1488 -3493 1488
rect -3459 -1488 -3453 1488
rect -3499 -1500 -3453 -1488
rect -3341 1488 -3295 1500
rect -3341 -1488 -3335 1488
rect -3301 -1488 -3295 1488
rect -3341 -1500 -3295 -1488
rect -3183 1488 -3137 1500
rect -3183 -1488 -3177 1488
rect -3143 -1488 -3137 1488
rect -3183 -1500 -3137 -1488
rect -3025 1488 -2979 1500
rect -3025 -1488 -3019 1488
rect -2985 -1488 -2979 1488
rect -3025 -1500 -2979 -1488
rect -2867 1488 -2821 1500
rect -2867 -1488 -2861 1488
rect -2827 -1488 -2821 1488
rect -2867 -1500 -2821 -1488
rect -2709 1488 -2663 1500
rect -2709 -1488 -2703 1488
rect -2669 -1488 -2663 1488
rect -2709 -1500 -2663 -1488
rect -2551 1488 -2505 1500
rect -2551 -1488 -2545 1488
rect -2511 -1488 -2505 1488
rect -2551 -1500 -2505 -1488
rect -2393 1488 -2347 1500
rect -2393 -1488 -2387 1488
rect -2353 -1488 -2347 1488
rect -2393 -1500 -2347 -1488
rect -2235 1488 -2189 1500
rect -2235 -1488 -2229 1488
rect -2195 -1488 -2189 1488
rect -2235 -1500 -2189 -1488
rect -2077 1488 -2031 1500
rect -2077 -1488 -2071 1488
rect -2037 -1488 -2031 1488
rect -2077 -1500 -2031 -1488
rect -1919 1488 -1873 1500
rect -1919 -1488 -1913 1488
rect -1879 -1488 -1873 1488
rect -1919 -1500 -1873 -1488
rect -1761 1488 -1715 1500
rect -1761 -1488 -1755 1488
rect -1721 -1488 -1715 1488
rect -1761 -1500 -1715 -1488
rect -1603 1488 -1557 1500
rect -1603 -1488 -1597 1488
rect -1563 -1488 -1557 1488
rect -1603 -1500 -1557 -1488
rect -1445 1488 -1399 1500
rect -1445 -1488 -1439 1488
rect -1405 -1488 -1399 1488
rect -1445 -1500 -1399 -1488
rect -1287 1488 -1241 1500
rect -1287 -1488 -1281 1488
rect -1247 -1488 -1241 1488
rect -1287 -1500 -1241 -1488
rect -1129 1488 -1083 1500
rect -1129 -1488 -1123 1488
rect -1089 -1488 -1083 1488
rect -1129 -1500 -1083 -1488
rect -971 1488 -925 1500
rect -971 -1488 -965 1488
rect -931 -1488 -925 1488
rect -971 -1500 -925 -1488
rect -813 1488 -767 1500
rect -813 -1488 -807 1488
rect -773 -1488 -767 1488
rect -813 -1500 -767 -1488
rect -655 1488 -609 1500
rect -655 -1488 -649 1488
rect -615 -1488 -609 1488
rect -655 -1500 -609 -1488
rect -497 1488 -451 1500
rect -497 -1488 -491 1488
rect -457 -1488 -451 1488
rect -497 -1500 -451 -1488
rect -339 1488 -293 1500
rect -339 -1488 -333 1488
rect -299 -1488 -293 1488
rect -339 -1500 -293 -1488
rect -181 1488 -135 1500
rect -181 -1488 -175 1488
rect -141 -1488 -135 1488
rect -181 -1500 -135 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 135 1488 181 1500
rect 135 -1488 141 1488
rect 175 -1488 181 1488
rect 135 -1500 181 -1488
rect 293 1488 339 1500
rect 293 -1488 299 1488
rect 333 -1488 339 1488
rect 293 -1500 339 -1488
rect 451 1488 497 1500
rect 451 -1488 457 1488
rect 491 -1488 497 1488
rect 451 -1500 497 -1488
rect 609 1488 655 1500
rect 609 -1488 615 1488
rect 649 -1488 655 1488
rect 609 -1500 655 -1488
rect 767 1488 813 1500
rect 767 -1488 773 1488
rect 807 -1488 813 1488
rect 767 -1500 813 -1488
rect 925 1488 971 1500
rect 925 -1488 931 1488
rect 965 -1488 971 1488
rect 925 -1500 971 -1488
rect 1083 1488 1129 1500
rect 1083 -1488 1089 1488
rect 1123 -1488 1129 1488
rect 1083 -1500 1129 -1488
rect 1241 1488 1287 1500
rect 1241 -1488 1247 1488
rect 1281 -1488 1287 1488
rect 1241 -1500 1287 -1488
rect 1399 1488 1445 1500
rect 1399 -1488 1405 1488
rect 1439 -1488 1445 1488
rect 1399 -1500 1445 -1488
rect 1557 1488 1603 1500
rect 1557 -1488 1563 1488
rect 1597 -1488 1603 1488
rect 1557 -1500 1603 -1488
rect 1715 1488 1761 1500
rect 1715 -1488 1721 1488
rect 1755 -1488 1761 1488
rect 1715 -1500 1761 -1488
rect 1873 1488 1919 1500
rect 1873 -1488 1879 1488
rect 1913 -1488 1919 1488
rect 1873 -1500 1919 -1488
rect 2031 1488 2077 1500
rect 2031 -1488 2037 1488
rect 2071 -1488 2077 1488
rect 2031 -1500 2077 -1488
rect 2189 1488 2235 1500
rect 2189 -1488 2195 1488
rect 2229 -1488 2235 1488
rect 2189 -1500 2235 -1488
rect 2347 1488 2393 1500
rect 2347 -1488 2353 1488
rect 2387 -1488 2393 1488
rect 2347 -1500 2393 -1488
rect 2505 1488 2551 1500
rect 2505 -1488 2511 1488
rect 2545 -1488 2551 1488
rect 2505 -1500 2551 -1488
rect 2663 1488 2709 1500
rect 2663 -1488 2669 1488
rect 2703 -1488 2709 1488
rect 2663 -1500 2709 -1488
rect 2821 1488 2867 1500
rect 2821 -1488 2827 1488
rect 2861 -1488 2867 1488
rect 2821 -1500 2867 -1488
rect 2979 1488 3025 1500
rect 2979 -1488 2985 1488
rect 3019 -1488 3025 1488
rect 2979 -1500 3025 -1488
rect 3137 1488 3183 1500
rect 3137 -1488 3143 1488
rect 3177 -1488 3183 1488
rect 3137 -1500 3183 -1488
rect 3295 1488 3341 1500
rect 3295 -1488 3301 1488
rect 3335 -1488 3341 1488
rect 3295 -1500 3341 -1488
rect 3453 1488 3499 1500
rect 3453 -1488 3459 1488
rect 3493 -1488 3499 1488
rect 3453 -1500 3499 -1488
rect 3611 1488 3657 1500
rect 3611 -1488 3617 1488
rect 3651 -1488 3657 1488
rect 3611 -1500 3657 -1488
rect 3769 1488 3815 1500
rect 3769 -1488 3775 1488
rect 3809 -1488 3815 1488
rect 3769 -1500 3815 -1488
rect 3927 1488 3973 1500
rect 3927 -1488 3933 1488
rect 3967 -1488 3973 1488
rect 3927 -1500 3973 -1488
rect 4085 1488 4131 1500
rect 4085 -1488 4091 1488
rect 4125 -1488 4131 1488
rect 4085 -1500 4131 -1488
rect 4243 1488 4289 1500
rect 4243 -1488 4249 1488
rect 4283 -1488 4289 1488
rect 4243 -1500 4289 -1488
rect 4401 1488 4447 1500
rect 4401 -1488 4407 1488
rect 4441 -1488 4447 1488
rect 4401 -1500 4447 -1488
rect 4559 1488 4605 1500
rect 4559 -1488 4565 1488
rect 4599 -1488 4605 1488
rect 4559 -1500 4605 -1488
rect 4717 1488 4763 1500
rect 4717 -1488 4723 1488
rect 4757 -1488 4763 1488
rect 4717 -1500 4763 -1488
rect 4875 1488 4921 1500
rect 4875 -1488 4881 1488
rect 4915 -1488 4921 1488
rect 4875 -1500 4921 -1488
rect 5033 1488 5079 1500
rect 5033 -1488 5039 1488
rect 5073 -1488 5079 1488
rect 5033 -1500 5079 -1488
rect 5191 1488 5237 1500
rect 5191 -1488 5197 1488
rect 5231 -1488 5237 1488
rect 5191 -1500 5237 -1488
rect 5349 1488 5395 1500
rect 5349 -1488 5355 1488
rect 5389 -1488 5395 1488
rect 5349 -1500 5395 -1488
rect 5507 1488 5553 1500
rect 5507 -1488 5513 1488
rect 5547 -1488 5553 1488
rect 5507 -1500 5553 -1488
rect 5665 1488 5711 1500
rect 5665 -1488 5671 1488
rect 5705 -1488 5711 1488
rect 5665 -1500 5711 -1488
rect 5823 1488 5869 1500
rect 5823 -1488 5829 1488
rect 5863 -1488 5869 1488
rect 5823 -1500 5869 -1488
rect 5981 1488 6027 1500
rect 5981 -1488 5987 1488
rect 6021 -1488 6027 1488
rect 5981 -1500 6027 -1488
rect 6139 1488 6185 1500
rect 6139 -1488 6145 1488
rect 6179 -1488 6185 1488
rect 6139 -1500 6185 -1488
rect 6297 1488 6343 1500
rect 6297 -1488 6303 1488
rect 6337 -1488 6343 1488
rect 6297 -1500 6343 -1488
rect 6455 1488 6501 1500
rect 6455 -1488 6461 1488
rect 6495 -1488 6501 1488
rect 6455 -1500 6501 -1488
rect 6613 1488 6659 1500
rect 6613 -1488 6619 1488
rect 6653 -1488 6659 1488
rect 6613 -1500 6659 -1488
rect 6771 1488 6817 1500
rect 6771 -1488 6777 1488
rect 6811 -1488 6817 1488
rect 6771 -1500 6817 -1488
rect 6929 1488 6975 1500
rect 6929 -1488 6935 1488
rect 6969 -1488 6975 1488
rect 6929 -1500 6975 -1488
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 15 l 0.5 m 1 nf 88 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
