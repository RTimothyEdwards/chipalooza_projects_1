magic
tech sky130A
magscale 1 2
timestamp 1713888873
<< pwell >>
rect -201 -90582 201 90582
<< psubdiff >>
rect -165 90512 -69 90546
rect 69 90512 165 90546
rect -165 90450 -131 90512
rect 131 90450 165 90512
rect -165 -90512 -131 -90450
rect 131 -90512 165 -90450
rect -165 -90546 -69 -90512
rect 69 -90546 165 -90512
<< psubdiffcont >>
rect -69 90512 69 90546
rect -165 -90450 -131 90450
rect 131 -90450 165 90450
rect -69 -90546 69 -90512
<< xpolycontact >>
rect -35 89984 35 90416
rect -35 -90416 35 -89984
<< ppolyres >>
rect -35 -89984 35 89984
<< locali >>
rect -165 90512 -69 90546
rect 69 90512 165 90546
rect -165 90450 -131 90512
rect 131 90450 165 90512
rect -165 -90512 -131 -90450
rect 131 -90512 165 -90450
rect -165 -90546 -69 -90512
rect 69 -90546 165 -90512
<< viali >>
rect -19 90001 19 90398
rect -19 -90398 19 -90001
<< metal1 >>
rect -25 90398 25 90410
rect -25 90001 -19 90398
rect 19 90001 25 90398
rect -25 89989 25 90001
rect -25 -90001 25 -89989
rect -25 -90398 -19 -90001
rect 19 -90398 25 -90001
rect -25 -90410 25 -90398
<< properties >>
string FIXED_BBOX -148 -90529 148 90529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 900.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 823.456k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
