magic
tech sky130A
magscale 1 2
timestamp 1714180253
<< psubdiff >>
rect 3348 5238 3808 5296
rect 3348 3328 3402 5238
rect 3750 3328 3808 5238
rect 3348 3288 3808 3328
<< psubdiffcont >>
rect 3402 3328 3750 5238
<< locali >>
rect 2942 6450 3028 6470
rect 2942 6126 2952 6450
rect 3016 6126 3028 6450
rect 2942 6112 3028 6126
rect 1184 5502 1430 5506
rect -1418 5456 -974 5470
rect -1418 5412 -1404 5456
rect -990 5412 -974 5456
rect -1418 5398 -974 5412
rect -908 5456 -464 5470
rect -908 5412 -890 5456
rect -486 5412 -464 5456
rect -908 5398 -464 5412
rect 1184 5374 1202 5502
rect 1410 5374 1430 5502
rect 1184 5366 1430 5374
rect -2291 5162 -2110 5297
rect -2291 4907 -2275 5162
rect -2124 4907 -2110 5162
rect 3340 5238 3794 5286
rect -1190 4992 -702 5096
rect 3340 5074 3402 5238
rect 886 4922 3402 5074
rect -2291 4890 -2110 4907
rect -4108 4734 -1552 4762
rect -4108 4642 -4090 4734
rect -1570 4642 -1552 4734
rect -4108 4636 -1552 4642
rect 160 4712 3046 4722
rect 160 4638 166 4712
rect 3036 4638 3046 4712
rect 160 4632 3046 4638
rect 3340 3328 3402 4922
rect 3750 3328 3794 5238
rect 3340 3294 3794 3328
<< viali >>
rect 2952 6126 3016 6450
rect -1404 5412 -990 5456
rect -890 5412 -486 5456
rect 1202 5374 1410 5502
rect -2275 4907 -2124 5162
rect -4090 4642 -1570 4734
rect 166 4638 3036 4712
<< metal1 >>
rect 896 6718 3020 6722
rect 558 6590 3020 6718
rect 558 6566 1128 6590
rect -1984 5802 410 6000
rect -2203 5480 -2085 5493
rect -2203 5386 -2192 5480
rect -2097 5386 -2085 5480
rect -2203 5375 -2085 5386
rect -2291 5162 -2110 5176
rect -2291 4907 -2275 5162
rect -2124 4907 -2110 5162
rect -2291 4890 -2110 4907
rect -1984 4780 -1518 5802
rect -1418 5456 -974 5470
rect -1418 5412 -1404 5456
rect -990 5412 -974 5456
rect -1418 5398 -974 5412
rect -908 5456 -250 5470
rect -908 5412 -890 5456
rect -486 5412 -250 5456
rect -908 5398 -250 5412
rect -4218 4734 -1518 4780
rect -1400 4848 -1328 5398
rect -1248 5118 -462 5176
rect -1248 4942 -1198 5118
rect -516 4942 -462 5118
rect -1248 4890 -462 4942
rect -1400 4776 -722 4848
rect -4218 4642 -4090 4734
rect -1570 4642 -1518 4734
rect -4218 4556 -1518 4642
rect -794 3498 -722 4776
rect -1150 3426 -722 3498
rect -322 3494 -250 5398
rect -66 4742 408 5802
rect 558 5182 816 6566
rect 2942 6460 3174 6470
rect 2942 6450 3090 6460
rect 2942 6126 2952 6450
rect 3016 6126 3090 6450
rect 2942 6122 3090 6126
rect 3158 6122 3174 6460
rect 2942 6112 3174 6122
rect 896 5760 3500 6004
rect 908 5694 2994 5710
rect 908 5642 948 5694
rect 2938 5642 2994 5694
rect 908 5630 2994 5642
rect 1184 5502 1430 5508
rect 1184 5374 1202 5502
rect 1410 5374 1430 5502
rect 1184 5366 1430 5374
rect 558 5176 1004 5182
rect 554 5082 3012 5176
rect 554 4958 928 5082
rect 2888 4958 3012 5082
rect 554 4890 3012 4958
rect 3218 4742 3500 5760
rect -66 4712 3500 4742
rect -66 4638 166 4712
rect 3036 4638 3500 4712
rect -66 4530 3500 4638
rect -66 4528 408 4530
rect -322 3422 139 3494
rect -664 2820 -406 2856
rect -1078 2544 234 2820
rect 3218 2780 3500 4530
rect -1078 2542 38 2544
rect -5530 2120 -4980 2360
rect 3930 2350 4452 2366
rect 3926 2120 4452 2350
rect -1258 1542 220 1750
rect -640 -288 -378 1542
rect 26 206 260 442
<< via1 >>
rect -2192 5386 -2097 5480
rect -2275 4907 -2124 5162
rect -1198 4942 -516 5118
rect 3090 6122 3158 6460
rect 948 5642 2938 5694
rect 1202 5374 1410 5502
rect 928 4958 2888 5082
<< metal2 >>
rect 3082 6460 3168 6470
rect 3082 6122 3090 6460
rect 3158 6122 3168 6460
rect -4360 5918 -4050 5924
rect -4360 5694 2994 5918
rect -4360 5642 948 5694
rect 2938 5642 2994 5694
rect -4360 5614 2994 5642
rect 1184 5502 1430 5508
rect -4370 5494 -4170 5498
rect 1184 5494 1202 5502
rect -4370 5480 1202 5494
rect -4370 5386 -2192 5480
rect -2097 5386 1202 5480
rect -4370 5374 1202 5386
rect 1410 5374 1430 5502
rect -4370 5372 1430 5374
rect -4370 5298 -4170 5372
rect 1184 5366 1430 5372
rect -4384 5162 2944 5176
rect -4384 4907 -2275 5162
rect -2124 5118 2944 5162
rect -2124 4942 -1198 5118
rect -516 5082 2944 5118
rect -516 4958 928 5082
rect 2888 4958 2944 5082
rect -516 4942 2944 4958
rect -2124 4907 2944 4942
rect -4384 4890 2944 4907
rect 3082 3530 3168 6122
rect 1632 3478 3168 3530
rect -5200 34 4112 438
use isolated_switch  isolated_switch_1
timestamp 1714078654
transform 1 0 -301 0 1 2911
box 301 -2911 4463 1830
use isolated_switch  isolated_switch_2
timestamp 1714078654
transform -1 0 -743 0 1 2911
box 301 -2911 4463 1830
use sky130_fd_pr__diode_pw2nd_05v5_HTFGEA  sky130_fd_pr__diode_pw2nd_05v5_HTFGEA_0  paramcells
timestamp 1714178384
transform 1 0 -2144 0 1 5433
box -186 -186 186 186
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform -1 0 -704 0 1 5089
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 896 0 1 5065
box -66 -43 2178 1671
<< labels >>
flabel metal1 -638 2556 -428 2832 0 FreeSans 560 0 0 0 avdd
port 4 nsew
flabel metal2 -970 156 -736 392 0 FreeSans 560 0 0 0 avss
port 5 nsew
flabel metal1 4234 2136 4436 2342 0 FreeSans 560 0 0 0 inA
port 6 nsew
flabel metal1 -604 -274 -400 -66 0 FreeSans 560 0 0 0 out
port 3 nsew
flabel metal1 -5504 2140 -5298 2338 0 FreeSans 560 0 0 0 inB
port 7 nsew
flabel metal2 -4360 5614 -4050 5924 0 FreeSans 560 0 0 0 dvdd
port 2 nsew
flabel metal2 -4384 4890 -4052 5176 0 FreeSans 560 0 0 0 dvss
port 0 nsew
flabel metal2 -4370 5298 -4170 5498 0 FreeSans 560 0 0 0 selA
port 1 nsew
<< end >>
