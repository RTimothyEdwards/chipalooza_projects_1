magic
tech sky130A
magscale 1 2
timestamp 1714090311
<< nwell >>
rect -362 -597 362 597
<< mvpmos >>
rect -100 -300 100 300
<< mvpdiff >>
rect -158 288 -100 300
rect -158 -288 -146 288
rect -112 -288 -100 288
rect -158 -300 -100 -288
rect 100 288 158 300
rect 100 -288 112 288
rect 146 -288 158 288
rect 100 -300 158 -288
<< mvpdiffc >>
rect -146 -288 -112 288
rect 112 -288 146 288
<< mvnsubdiff >>
rect -296 519 296 531
rect -296 485 -184 519
rect 184 485 296 519
rect -296 473 296 485
rect -296 423 -238 473
rect -296 -423 -284 423
rect -250 -423 -238 423
rect 238 423 296 473
rect -296 -473 -238 -423
rect 238 -423 250 423
rect 284 -423 296 423
rect 238 -473 296 -423
rect -296 -485 296 -473
rect -296 -519 -184 -485
rect 184 -519 296 -485
rect -296 -531 296 -519
<< mvnsubdiffcont >>
rect -184 485 184 519
rect -284 -423 -250 423
rect 250 -423 284 423
rect -184 -519 184 -485
<< poly >>
rect -100 381 100 397
rect -100 347 -84 381
rect 84 347 100 381
rect -100 300 100 347
rect -100 -347 100 -300
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -397 100 -381
<< polycont >>
rect -84 347 84 381
rect -84 -381 84 -347
<< locali >>
rect -284 485 -184 519
rect 184 485 284 519
rect -284 423 -250 485
rect 250 423 284 485
rect -100 347 -84 381
rect 84 347 100 381
rect -146 288 -112 304
rect -146 -304 -112 -288
rect 112 288 146 304
rect 112 -304 146 -288
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -284 -485 -250 -423
rect 250 -485 284 -423
rect -284 -519 -184 -485
rect 184 -519 284 -485
<< viali >>
rect -284 -388 -250 388
rect -84 347 84 381
rect -146 -288 -112 288
rect 112 -288 146 288
rect -84 -381 84 -347
rect 250 -388 284 388
<< metal1 >>
rect -290 388 -244 400
rect -290 -388 -284 388
rect -250 -388 -244 388
rect 244 388 290 400
rect -96 381 96 387
rect -96 347 -84 381
rect 84 347 96 381
rect -96 341 96 347
rect -152 288 -106 300
rect -152 -288 -146 288
rect -112 -288 -106 288
rect -152 -300 -106 -288
rect 106 288 152 300
rect 106 -288 112 288
rect 146 -288 152 288
rect 106 -300 152 -288
rect -96 -347 96 -341
rect -96 -381 -84 -347
rect 84 -381 96 -347
rect -96 -387 96 -381
rect -290 -400 -244 -388
rect 244 -388 250 388
rect 284 -388 290 388
rect 244 -400 290 -388
<< properties >>
string FIXED_BBOX -263 -502 263 502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 80 viagl 80 viagt 0
<< end >>
