magic
tech sky130A
magscale 1 2
timestamp 1713984708
<< metal1 >>
rect -20400 3360 -9499 49600
rect -85199 -10677 -23576 -9757
rect -85199 -28067 -79389 -10677
rect -78189 -28067 -67389 -10677
rect -66189 -28067 -55389 -10677
rect -54189 -28067 -43389 -10677
rect -42189 -28067 -31389 -10677
rect -30189 -28067 -23576 -10677
rect -85199 -30024 -23576 -28067
rect -21510 -29400 -21500 -13300
rect -21160 -29400 -21150 -13300
rect -15450 -29400 -15440 -13300
rect -15100 -29400 -15090 -13300
rect -85209 -32280 -85199 -30024
rect -23576 -32280 -23566 -30024
<< via1 >>
rect -21500 -29400 -21160 -13300
rect -15440 -29400 -15100 -13300
rect -85199 -32280 -23576 -30024
<< metal2 >>
rect -20400 3360 -9499 49600
rect -22348 422 -16669 423
rect -22350 -50 -16669 422
rect -22822 -1386 -16669 -50
rect -22342 -1388 -16669 -1386
rect -85199 -10677 -23576 -9757
rect -85199 -28067 -79389 -10677
rect -78189 -28067 -67389 -10677
rect -66189 -28067 -55389 -10677
rect -54189 -28067 -43389 -10677
rect -42189 -28067 -31389 -10677
rect -30189 -28067 -23576 -10677
rect -85199 -30024 -23576 -28067
rect -21900 -13290 -21160 -13280
rect -18340 -13418 -16669 -1388
rect -15440 -13300 -14700 -13290
rect -21900 -29420 -21160 -29410
rect -16566 -29414 -16506 -28852
rect -85199 -32290 -23576 -32280
rect -16682 -29474 -16506 -29414
rect -16462 -29415 -16402 -28852
rect -15440 -29410 -14700 -29400
rect -16682 -44204 -16622 -29474
rect -16462 -29475 -16262 -29415
rect -16322 -44204 -16262 -29475
<< via2 >>
rect -21900 -13300 -21160 -13290
rect -21900 -29400 -21500 -13300
rect -21500 -29400 -21160 -13300
rect -21900 -29410 -21160 -29400
rect -85199 -32280 -23576 -30024
rect -15440 -29400 -15100 -13300
rect -15100 -29400 -14700 -13300
<< metal3 >>
rect -89200 -4000 -79200 66802
rect -75200 56800 -9502 66800
rect -18400 43364 -9502 56800
rect -18400 3411 -9500 43364
rect -20400 1520 -9500 3411
rect -89200 -4576 -22388 -4000
rect -89200 -11276 -21135 -4576
rect -89200 -12561 -82816 -11276
rect -25932 -12561 -21135 -11276
rect -89200 -13290 -21135 -12561
rect -89200 -18044 -21900 -13290
rect -89200 -19329 -82559 -18044
rect -25675 -19329 -21900 -18044
rect -89200 -24000 -21900 -19329
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11471 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11471 -13300
rect -85209 -30024 -23566 -30019
rect -15464 -30024 -11471 -29400
rect -87200 -32280 -85199 -30024
rect -23576 -32280 -11471 -30024
rect -87200 -37148 -11471 -32280
rect -87200 -38433 -79646 -37148
rect -22762 -38433 -11471 -37148
rect -87200 -44000 -11471 -38433
<< via3 >>
rect -21900 -29410 -21160 -13290
rect -15440 -29400 -14700 -13300
rect -85199 -32280 -23576 -30024
<< metal4 >>
rect -89200 -4000 -79200 66802
rect -75200 56800 -9502 66800
rect -18400 43364 -9502 56800
rect -18400 3411 -9500 43364
rect -20400 1520 -9500 3411
rect -89200 -4576 -22388 -4000
rect -89200 -11276 -21135 -4576
rect -89200 -12561 -82816 -11276
rect -25932 -12561 -21135 -11276
rect -89200 -13290 -21135 -12561
rect -89200 -18044 -21900 -13290
rect -89200 -19329 -82559 -18044
rect -25675 -19329 -21900 -18044
rect -89200 -24000 -21900 -19329
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11471 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11471 -13300
rect -85200 -30024 -23575 -30023
rect -15464 -30024 -11471 -29400
rect -87200 -32280 -85199 -30024
rect -23576 -32280 -11471 -30024
rect -87200 -37148 -11471 -32280
rect -87200 -38433 -79646 -37148
rect -22762 -38433 -11471 -37148
rect -87200 -44000 -11471 -38433
<< via4 >>
rect -21900 -29410 -21160 -13290
rect -15440 -29400 -14700 -13300
rect -85199 -32280 -23576 -30024
<< metal5 >>
rect -89200 -4000 -79200 66802
rect -75200 56800 -9502 66800
rect -18400 43364 -9502 56800
rect -18400 3411 -9500 43364
rect -20400 1520 -9500 3411
rect -89200 -4576 -22388 -4000
rect -89200 -11276 -21135 -4576
rect -89200 -12561 -82816 -11276
rect -25932 -12561 -21135 -11276
rect -89200 -13290 -21135 -12561
rect -89200 -18044 -21900 -13290
rect -89200 -19329 -82559 -18044
rect -25675 -19329 -21900 -18044
rect -89200 -24000 -21900 -19329
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11471 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11471 -13300
rect -21924 -29434 -21136 -29433
rect -85223 -30024 -23552 -30000
rect -15464 -30024 -11471 -29400
rect -87200 -32280 -85199 -30024
rect -23576 -32280 -11471 -30024
rect -87200 -37148 -11471 -32280
rect -87200 -38433 -79646 -37148
rect -22762 -38433 -11471 -37148
rect -87200 -44000 -11471 -38433
use gate_drive  gate_drive_0
timestamp 1624430562
transform 0 -1 -17500 1 0 -20900
box -8500 -2400 7600 4000
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1624430562
transform -1 0 -22400 0 1 0
box -10800 -10800 63600 63600
<< labels >>
flabel metal5 -89200 66679 -79200 66802 5 FreeSans 8000 0 0 0 vdd_pwr
port 9 s
flabel metal5 -87200 -44000 -87179 -30024 1 FreeSans 8000 0 0 0 vss
port 10 n
flabel metal2 -16322 -44204 -16262 -44203 1 FreeSans 400 0 0 0 p_in_n
port 4 n
flabel metal2 -16682 -44204 -16622 -44203 1 FreeSans 400 0 0 0 p_in
port 3 n
flabel metal5 -75200 65820 -9502 66800 1 FreeSans 8000 0 0 0 sw_node
port 7 n
<< end >>
