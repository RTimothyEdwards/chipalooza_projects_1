magic
tech sky130A
magscale 1 2
timestamp 1713995538
<< pwell >>
rect -453 -5169 -383 -4737
rect 15100 -5541 15188 -5406
<< locali >>
rect 35266 -3135 35328 -2897
<< metal1 >>
rect -583 1818 12861 1829
rect -583 1766 -550 1818
rect 12825 1766 12861 1818
rect -583 1754 12861 1766
rect -583 1431 -383 1663
rect -902 1231 -383 1431
rect -287 1231 -51 1663
rect 45 1231 281 1663
rect 377 1231 613 1663
rect 709 1231 945 1663
rect 1041 1231 1277 1663
rect 1373 1231 1609 1663
rect 1705 1231 1941 1663
rect 2037 1231 2273 1663
rect 2369 1231 2605 1663
rect 2701 1231 2937 1663
rect 3033 1231 3269 1663
rect 3365 1231 3601 1663
rect 3697 1231 3933 1663
rect 4029 1231 4265 1663
rect 4361 1231 4597 1663
rect 4693 1231 4929 1663
rect 5025 1231 5261 1663
rect 5357 1231 5593 1663
rect 5689 1231 5925 1663
rect 6021 1231 6257 1663
rect 6353 1231 6589 1663
rect 6685 1231 6921 1663
rect 7017 1231 7253 1663
rect 7349 1231 7585 1663
rect -589 -4869 -537 1069
rect 7681 577 7917 1663
rect 8013 1231 8249 1663
rect 8345 1231 8581 1663
rect 8677 1231 8913 1663
rect 9009 1231 9245 1663
rect 9341 1231 9577 1663
rect 9673 1231 9909 1663
rect 10005 1231 10241 1663
rect 10337 1231 10573 1663
rect 10669 1231 10905 1663
rect 11001 1231 11237 1663
rect 11333 1231 11569 1663
rect 11665 1231 11901 1663
rect 11997 1231 12233 1663
rect 12329 1231 12565 1663
rect 12660 1371 12861 1663
rect 12660 1231 13108 1371
rect 7681 328 7917 343
rect 12821 -1873 12873 -1859
rect 12821 -2125 12873 -2111
rect 12968 -3739 13108 1231
rect 46289 -427 46357 -318
rect 46139 -661 46289 -459
rect 46139 -705 46357 -661
rect 14752 -3228 14814 -2882
rect 15278 -3228 15340 -2882
rect 15804 -3228 15866 -2882
rect 16330 -3228 16392 -2882
rect 16856 -3228 16918 -2882
rect 17382 -3228 17444 -2882
rect 17908 -3228 17970 -2882
rect 18434 -3228 18496 -2882
rect 18960 -3228 19022 -2882
rect 19486 -3228 19548 -2882
rect 20012 -3228 20074 -2882
rect 20538 -3228 20600 -2882
rect 21064 -3228 21126 -2882
rect 21590 -3228 21652 -2882
rect 22116 -3228 22178 -2882
rect 22642 -3228 22704 -2882
rect 23168 -3228 23230 -2882
rect 23694 -3228 23756 -2882
rect 24220 -3228 24282 -2882
rect 24746 -3228 24808 -2882
rect 25272 -3228 25334 -2882
rect 25798 -3228 25860 -2882
rect 26324 -3228 26386 -2882
rect 26850 -3228 26912 -2882
rect 27376 -3228 27438 -2882
rect 27902 -3228 27964 -2882
rect 28428 -3228 28490 -2882
rect 28954 -3228 29016 -2882
rect 29480 -3228 29542 -2882
rect 30006 -3228 30068 -2882
rect 30532 -3228 30594 -2882
rect 31058 -3228 31120 -2882
rect 31584 -3228 31646 -2882
rect 32110 -3228 32172 -2882
rect 32636 -3228 32698 -2882
rect 33162 -3228 33224 -2882
rect 33688 -3228 33750 -2882
rect 34214 -3228 34276 -2882
rect 34740 -3228 34802 -2882
rect 35266 -3228 35328 -2882
rect 35792 -2897 35854 -2882
rect 35792 -3228 35854 -3135
rect 36318 -2897 36380 -2882
rect 36318 -3228 36380 -3135
rect 36844 -2897 36906 -2882
rect 36844 -3228 36906 -3135
rect 37370 -2897 37432 -2882
rect 37370 -3228 37432 -3135
rect 37896 -2897 37958 -2882
rect 37896 -3228 37958 -3135
rect 38422 -2897 38484 -2882
rect 38422 -3228 38484 -3135
rect 38948 -2897 39010 -2882
rect 38948 -3228 39010 -3135
rect 39474 -2897 39536 -2882
rect 39474 -3228 39536 -3135
rect 40000 -2897 40062 -2882
rect 40000 -3228 40062 -3135
rect 40526 -2897 40588 -2882
rect 40526 -3228 40588 -3135
rect 41052 -2897 41114 -2882
rect 41052 -3228 41114 -3135
rect 41578 -2897 41640 -2882
rect 41578 -3228 41640 -3135
rect 42104 -2897 42166 -2882
rect 42104 -3228 42166 -3135
rect 42630 -2897 42692 -2882
rect 42630 -3228 42692 -3135
rect 43156 -2897 43218 -2882
rect 43156 -3228 43218 -3135
rect 43682 -2897 43744 -2882
rect 43682 -3228 43744 -3135
rect 44208 -2897 44270 -2882
rect 44208 -3228 44270 -3135
rect 44734 -2897 44796 -2882
rect 44734 -3228 44796 -3135
rect 45260 -2897 45322 -2882
rect 45260 -3228 45322 -3135
rect 45786 -2897 45848 -2882
rect 45786 -3228 45848 -3135
rect 14418 -4194 14482 -3871
rect 14944 -4194 15008 -3871
rect 15470 -4194 15534 -3871
rect 15996 -4194 16060 -3871
rect 16522 -4194 16586 -3871
rect 17048 -4194 17112 -3871
rect 17574 -4194 17638 -3871
rect 18100 -4194 18164 -3871
rect 18626 -4194 18690 -3871
rect 19152 -4194 19216 -3871
rect 19678 -4194 19742 -3871
rect 20204 -4194 20268 -3871
rect 20730 -4194 20794 -3871
rect 21256 -4194 21320 -3871
rect 21782 -4194 21846 -3871
rect 22308 -4194 22372 -3871
rect 22834 -4194 22898 -3871
rect 23360 -4194 23424 -3871
rect 23886 -4194 23950 -3871
rect 24412 -4194 24476 -3871
rect 24938 -4194 25002 -3871
rect 25464 -4194 25528 -3871
rect 25990 -4194 26054 -3871
rect 26516 -4194 26580 -3871
rect 27042 -4194 27106 -3871
rect 27568 -4194 27632 -3871
rect 28094 -4194 28158 -3871
rect 28620 -4194 28684 -3871
rect 29146 -4194 29210 -3871
rect 29672 -4194 29736 -3871
rect 30198 -4194 30262 -3871
rect 30724 -4194 30788 -3871
rect 31250 -4194 31314 -3871
rect 31776 -4194 31840 -3871
rect 32302 -4194 32366 -3871
rect 32828 -4194 32892 -3871
rect 33354 -4194 33418 -3871
rect 33880 -4194 33944 -3871
rect 34406 -4194 34470 -3871
rect 34932 -4194 34996 -3871
rect 35458 -4194 35522 -3871
rect 35984 -3881 36048 -3871
rect 35984 -4194 36048 -4119
rect 36510 -3881 36574 -3871
rect 36510 -4194 36574 -4119
rect 37036 -3881 37100 -3871
rect 37036 -4194 37100 -4119
rect 37562 -3881 37626 -3871
rect 37562 -4194 37626 -4119
rect 38088 -3881 38152 -3871
rect 38088 -4194 38152 -4119
rect 38614 -3881 38678 -3871
rect 38614 -4194 38678 -4119
rect 39140 -3881 39204 -3871
rect 39140 -4194 39204 -4119
rect 39666 -3881 39730 -3871
rect 39666 -4194 39730 -4119
rect 40192 -3881 40256 -3871
rect 40192 -4194 40256 -4119
rect 40718 -3881 40782 -3871
rect 40718 -4194 40782 -4119
rect 41244 -3881 41308 -3871
rect 41244 -4194 41308 -4119
rect 41770 -3881 41834 -3871
rect 41770 -4194 41834 -4119
rect 42296 -3881 42360 -3871
rect 42296 -4194 42360 -4119
rect 42822 -3881 42886 -3871
rect 42822 -4194 42886 -4119
rect 43348 -3881 43412 -3871
rect 43348 -4194 43412 -4119
rect 43874 -3881 43938 -3871
rect 43874 -4194 43938 -4119
rect 44400 -3881 44464 -3871
rect 44400 -4194 44464 -4119
rect 44926 -3881 44990 -3871
rect 44926 -4194 44990 -4119
rect 45452 -3881 45516 -3871
rect 45452 -4194 45516 -4119
rect 12968 -4262 13108 -4225
rect -589 -5305 -537 -5107
rect -453 -5169 -217 -4737
rect -121 -5169 115 -4737
rect 211 -5169 447 -4737
rect 543 -5169 779 -4737
rect 875 -5169 1111 -4737
rect 1207 -5169 1443 -4737
rect 1539 -5169 1775 -4737
rect 1871 -5169 2107 -4737
rect 2203 -5169 2439 -4737
rect 2535 -5169 2771 -4737
rect 2867 -5169 3103 -4737
rect 3199 -5169 3435 -4737
rect 3531 -5169 3767 -4737
rect 3863 -5169 4099 -4737
rect 4195 -5169 4431 -4737
rect 4527 -5169 4763 -4737
rect 4859 -5169 5095 -4737
rect 5191 -5169 5427 -4737
rect 5523 -5169 5759 -4737
rect 5855 -5169 6091 -4737
rect 6187 -5169 6423 -4737
rect 6519 -5169 6755 -4737
rect 6851 -5169 7087 -4737
rect 7183 -5169 7419 -4737
rect 7515 -5169 7751 -4737
rect 7847 -5169 8083 -4737
rect 8179 -5169 8415 -4737
rect 8511 -5169 8747 -4737
rect 8843 -5169 9079 -4737
rect 9175 -5169 9411 -4737
rect 9507 -5169 9743 -4737
rect 9839 -5169 10075 -4737
rect 10171 -5169 10407 -4737
rect 10503 -5169 10739 -4737
rect 10835 -5169 11071 -4737
rect 11167 -5169 11403 -4737
rect 11499 -5169 11735 -4737
rect 11831 -5169 12067 -4737
rect 12163 -5169 12399 -4737
rect 12495 -5169 12731 -4737
rect 12821 -5305 12867 -4575
rect 15110 -5532 15164 -5316
rect 15636 -5532 15690 -5316
rect 16162 -5532 16216 -5316
rect 16688 -5532 16742 -5316
rect 17214 -5532 17268 -5316
rect 17740 -5532 17794 -5316
rect 18266 -5532 18320 -5316
rect 18792 -5532 18846 -5316
rect 19318 -5532 19372 -5316
rect 19844 -5532 19898 -5316
rect 20370 -5532 20424 -5316
rect 20896 -5532 20950 -5316
rect 21422 -5532 21476 -5316
rect 21948 -5532 22002 -5316
rect 22474 -5532 22528 -5316
rect 23000 -5532 23054 -5316
rect 23526 -5532 23580 -5316
rect 24052 -5532 24106 -5316
rect 24578 -5532 24632 -5316
rect 25104 -5532 25158 -5316
rect 25630 -5532 25684 -5316
rect 26156 -5532 26210 -5316
rect 26682 -5532 26736 -5316
rect 27208 -5532 27262 -5316
rect 27734 -5532 27788 -5316
rect 28260 -5532 28314 -5316
rect 28786 -5532 28840 -5316
rect 29312 -5532 29366 -5316
rect 29838 -5532 29892 -5316
rect 30364 -5532 30418 -5316
rect 30890 -5532 30944 -5316
rect 31416 -5532 31470 -5316
rect 31942 -5532 31996 -5316
rect 32468 -5532 32522 -5316
rect 32994 -5532 33048 -5316
rect 33520 -5532 33574 -5316
rect 34046 -5532 34100 -5316
rect 34572 -5532 34626 -5316
rect 35098 -5532 35152 -5316
rect 35624 -5532 35678 -5316
rect 36150 -5532 36204 -5504
rect 36676 -5532 36730 -5504
rect 37202 -5532 37256 -5504
rect 37728 -5532 37782 -5504
rect 38254 -5532 38308 -5504
rect 38780 -5532 38834 -5504
rect 39306 -5532 39360 -5504
rect 39832 -5532 39886 -5504
rect 40358 -5532 40412 -5504
rect 40884 -5532 40938 -5504
rect 41410 -5532 41464 -5504
rect 41936 -5532 41990 -5504
rect 42462 -5532 42516 -5504
rect 42988 -5532 43042 -5504
rect 43514 -5532 43568 -5504
rect 44040 -5532 44094 -5504
rect 44566 -5532 44620 -5504
rect 45092 -5532 45146 -5504
rect 45618 -5532 45672 -5504
rect 46144 -5532 46198 -5504
<< via1 >>
rect 46143 2384 46197 2616
rect -550 1766 12825 1818
rect 7681 343 7917 577
rect 12821 -2111 12873 -1873
rect 45984 677 46053 1236
rect 46289 -661 46357 -427
rect 35792 -3135 35854 -2897
rect 36318 -3135 36380 -2897
rect 36844 -3135 36906 -2897
rect 37370 -3135 37432 -2897
rect 37896 -3135 37958 -2897
rect 38422 -3135 38484 -2897
rect 38948 -3135 39010 -2897
rect 39474 -3135 39536 -2897
rect 40000 -3135 40062 -2897
rect 40526 -3135 40588 -2897
rect 41052 -3135 41114 -2897
rect 41578 -3135 41640 -2897
rect 42104 -3135 42166 -2897
rect 42630 -3135 42692 -2897
rect 43156 -3135 43218 -2897
rect 43682 -3135 43744 -2897
rect 44208 -3135 44270 -2897
rect 44734 -3135 44796 -2897
rect 45260 -3135 45322 -2897
rect 45786 -3135 45848 -2897
rect 12968 -4225 13108 -3739
rect 35984 -4119 36048 -3881
rect 36510 -4119 36574 -3881
rect 37036 -4119 37100 -3881
rect 37562 -4119 37626 -3881
rect 38088 -4119 38152 -3881
rect 38614 -4119 38678 -3881
rect 39140 -4119 39204 -3881
rect 39666 -4119 39730 -3881
rect 40192 -4119 40256 -3881
rect 40718 -4119 40782 -3881
rect 41244 -4119 41308 -3881
rect 41770 -4119 41834 -3881
rect 42296 -4119 42360 -3881
rect 42822 -4119 42886 -3881
rect 43348 -4119 43412 -3881
rect 43874 -4119 43938 -3881
rect 44400 -4119 44464 -3881
rect 44926 -4119 44990 -3881
rect 45452 -4119 45516 -3881
rect -589 -5107 -537 -4869
rect 45978 -4774 46066 -4207
rect 36150 -5504 36204 -5316
rect 36676 -5504 36730 -5316
rect 37202 -5504 37256 -5316
rect 37728 -5504 37782 -5316
rect 38254 -5504 38308 -5316
rect 38780 -5504 38834 -5316
rect 39306 -5504 39360 -5316
rect 39832 -5504 39886 -5316
rect 40358 -5504 40412 -5316
rect 40884 -5504 40938 -5316
rect 41410 -5504 41464 -5316
rect 41936 -5504 41990 -5316
rect 42462 -5504 42516 -5316
rect 42988 -5504 43042 -5316
rect 43514 -5504 43568 -5316
rect 44040 -5504 44094 -5316
rect 44566 -5504 44620 -5316
rect 45092 -5504 45146 -5316
rect 45618 -5504 45672 -5316
rect 46144 -5504 46198 -5316
<< metal2 >>
rect 46082 2616 46242 2884
rect 13336 2382 13479 2614
rect 13685 2382 13944 2614
rect 14389 2382 45815 2614
rect 45901 2382 45910 2614
rect 46082 2384 46143 2616
rect 46197 2384 46242 2616
rect 13522 2075 13815 2307
rect 14021 2075 14120 2307
rect 14389 2075 45817 2307
rect 45903 2075 45914 2307
rect 46082 2065 46242 2384
rect 46279 2382 46289 2614
rect 46375 2382 54509 2614
rect 54836 2382 119979 2614
rect 120121 2382 164959 2614
rect 165286 2382 225185 2614
rect 225320 2382 228619 2614
rect 228946 2382 231498 2614
rect 231626 2382 233879 2614
rect 234206 2382 235691 2614
rect 235834 2382 237049 2614
rect 237376 2382 237806 2614
rect 237938 2382 239141 2614
rect 239468 2382 239910 2614
rect 240042 2382 241233 2614
rect 241560 2382 242014 2614
rect 242146 2382 242785 2614
rect 243112 2382 243126 2614
rect 243198 2382 243214 2614
rect 243386 2382 243420 2614
rect 243723 2382 243895 2614
rect 244112 2382 244330 2614
rect 46278 2075 46289 2307
rect 46375 2075 53614 2307
rect 53799 2075 119979 2307
rect 120121 2075 164064 2307
rect 164249 2075 225185 2307
rect 225320 2075 227724 2307
rect 227909 2075 231498 2307
rect 231626 2075 232984 2307
rect 233169 2075 235691 2307
rect 235834 2075 236154 2307
rect 236339 2075 237806 2307
rect 237938 2075 238246 2307
rect 238431 2075 239910 2307
rect 240042 2075 240338 2307
rect 240523 2075 242014 2307
rect 242146 2075 242430 2307
rect 242615 2075 243075 2307
rect 243198 2075 243556 2307
rect 243741 2075 243766 2307
rect 243910 2075 244239 2307
rect 244414 2075 244509 2307
rect -900 1818 12943 1912
rect -900 1766 -550 1818
rect 12825 1766 12943 1818
rect -900 1674 12943 1766
rect 13184 1674 14481 1912
rect -671 1343 13193 1577
rect 244825 1343 244872 1577
rect 245127 1343 245156 1577
rect 45984 1236 46053 1245
rect 45984 668 46053 677
rect -656 343 7681 577
rect 7917 343 14323 577
rect 12960 342 13191 343
rect 244825 -1715 244871 -1481
rect 245126 -1715 245155 -1481
rect 12811 -2111 12821 -1873
rect 12873 -2111 12944 -1873
rect 13185 -1892 14284 -1873
rect 13185 -1976 13323 -1892
rect 13185 -2111 14284 -1976
rect 14752 -3135 14814 -2897
rect 15278 -3135 15340 -2897
rect 15804 -3135 15866 -2897
rect 16330 -3135 16392 -2897
rect 16856 -3135 16918 -2897
rect 17382 -3135 17444 -2897
rect 17908 -3135 17970 -2897
rect 18434 -3135 18496 -2897
rect 18960 -3135 19022 -2897
rect 19486 -3135 19548 -2897
rect 20012 -3135 20074 -2897
rect 20538 -3135 20600 -2897
rect 21064 -3135 21126 -2897
rect 21590 -3135 21652 -2897
rect 22116 -3135 22178 -2897
rect 22642 -3135 22704 -2897
rect 23168 -3135 23230 -2897
rect 23694 -3135 23756 -2897
rect 24220 -3135 24282 -2897
rect 24746 -3135 24808 -2897
rect 25272 -3135 25334 -2897
rect 25798 -3135 25860 -2897
rect 26324 -3135 26386 -2897
rect 26850 -3135 26912 -2897
rect 27376 -3135 27438 -2897
rect 27902 -3135 27964 -2897
rect 28428 -3135 28490 -2897
rect 28954 -3135 29016 -2897
rect 29480 -3135 29542 -2897
rect 30006 -3135 30068 -2897
rect 30532 -3135 30594 -2897
rect 31058 -3135 31120 -2897
rect 31584 -3135 31646 -2897
rect 32110 -3135 32172 -2897
rect 32636 -3135 32698 -2897
rect 33162 -3135 33224 -2897
rect 33688 -3135 33750 -2897
rect 34214 -3135 34276 -2897
rect 34740 -3135 34802 -2897
rect 12956 -4225 12968 -3739
rect 13108 -3881 13119 -3739
rect 13108 -4119 35984 -3881
rect 36048 -4119 36510 -3881
rect 36574 -4119 37036 -3881
rect 37100 -4119 37562 -3881
rect 37626 -4119 38088 -3881
rect 38152 -4119 38614 -3881
rect 38678 -4119 39140 -3881
rect 39204 -4119 39666 -3881
rect 39730 -4119 40192 -3881
rect 40256 -4119 40718 -3881
rect 40782 -4119 41244 -3881
rect 41308 -4119 41770 -3881
rect 41834 -4119 42296 -3881
rect 42360 -4119 42822 -3881
rect 42886 -4119 43348 -3881
rect 43412 -4119 43874 -3881
rect 43938 -4119 44400 -3881
rect 44464 -4119 44926 -3881
rect 44990 -4119 45452 -3881
rect 45516 -4119 244806 -3881
rect 13108 -4225 13119 -4119
rect 12956 -4226 13119 -4225
rect 45978 -4207 46066 -4198
rect 45978 -4783 46066 -4774
rect -612 -5107 -589 -4869
rect -537 -5107 12944 -4869
rect 13185 -5107 14284 -4869
rect 12915 -5504 12944 -5316
rect 13070 -5504 14125 -5316
rect 14193 -5504 23221 -5316
rect 23406 -5504 35180 -5316
rect 35244 -5504 36150 -5316
rect 36204 -5504 36676 -5316
rect 36730 -5504 37202 -5316
rect 37256 -5504 37728 -5316
rect 37782 -5504 38254 -5316
rect 38308 -5504 38780 -5316
rect 38834 -5504 39306 -5316
rect 39360 -5504 39832 -5316
rect 39886 -5504 40358 -5316
rect 40412 -5504 40884 -5316
rect 40938 -5504 41410 -5316
rect 41464 -5504 41936 -5316
rect 41990 -5504 42462 -5316
rect 42516 -5504 42988 -5316
rect 43042 -5504 43514 -5316
rect 43568 -5504 44040 -5316
rect 44094 -5504 44566 -5316
rect 44620 -5504 45092 -5316
rect 45146 -5504 45618 -5316
rect 45672 -5504 46144 -5316
rect 46198 -5504 46372 -5316
rect 46661 -5504 69421 -5316
rect 69606 -5504 98806 -5316
rect 99244 -5504 122021 -5316
rect 122206 -5504 151424 -5316
rect 151834 -5504 174621 -5316
rect 174806 -5504 204020 -5316
rect 204444 -5504 227221 -5316
rect 227406 -5504 243456 -5316
rect 243907 -5504 244285 -5316
rect 244402 -5504 244517 -5316
rect 13355 -5760 13541 -5572
rect 13741 -5760 13965 -5572
rect 14412 -5760 24116 -5572
rect 24443 -5760 35012 -5572
rect 35244 -5590 35344 -5504
rect 35144 -5790 35344 -5590
rect 35430 -5760 45532 -5572
rect 45956 -5760 46048 -5572
rect 46498 -5760 70316 -5572
rect 70643 -5760 98652 -5572
rect 99090 -5760 122916 -5572
rect 123243 -5760 151268 -5572
rect 151678 -5760 175516 -5572
rect 175843 -5760 203868 -5572
rect 204292 -5760 228116 -5572
rect 228443 -5760 243298 -5572
rect 243742 -5760 243897 -5572
rect 244079 -5760 244352 -5572
<< via2 >>
rect 13479 2382 13685 2614
rect 45815 2382 45901 2614
rect 13815 2075 14021 2307
rect 45817 2075 45903 2307
rect 46289 2382 46375 2614
rect 54509 2382 54836 2614
rect 164959 2382 165286 2614
rect 228619 2382 228946 2614
rect 233879 2382 234206 2614
rect 237049 2382 237376 2614
rect 239141 2382 239468 2614
rect 241233 2382 241560 2614
rect 242785 2382 243112 2614
rect 243214 2382 243386 2614
rect 243895 2382 244112 2614
rect 46289 2075 46375 2307
rect 53614 2075 53799 2307
rect 164064 2075 164249 2307
rect 227724 2075 227909 2307
rect 232984 2075 233169 2307
rect 236154 2075 236339 2307
rect 238246 2075 238431 2307
rect 240338 2075 240523 2307
rect 242430 2075 242615 2307
rect 243556 2075 243741 2307
rect 244239 2075 244414 2307
rect 12943 1674 13184 1912
rect 244872 1343 245127 1577
rect 45984 677 46053 1236
rect 13322 -1699 45823 -1615
rect 46232 -1699 244671 -1615
rect 244871 -1715 245126 -1481
rect 12944 -2111 13185 -1873
rect 13323 -1976 45824 -1892
rect 46233 -1974 244672 -1890
rect 45978 -4774 46066 -4207
rect 12944 -5107 13185 -4869
rect 12944 -5504 13070 -5316
rect 23221 -5504 23406 -5316
rect 69421 -5504 69606 -5316
rect 122021 -5504 122206 -5316
rect 174621 -5504 174806 -5316
rect 227221 -5504 227406 -5316
rect 244285 -5504 244402 -5316
rect 13541 -5760 13741 -5572
rect 24116 -5760 24443 -5572
rect 70316 -5760 70643 -5572
rect 122916 -5760 123243 -5572
rect 175516 -5760 175843 -5572
rect 228116 -5760 228443 -5572
rect 243897 -5760 244079 -5572
<< metal3 >>
rect 13467 2614 13696 2928
rect 13467 2382 13479 2614
rect 13685 2382 13696 2614
rect 13467 2369 13696 2382
rect 13803 2307 14032 2928
rect 45809 2614 46383 2622
rect 45809 2382 45815 2614
rect 45901 2382 46289 2614
rect 46375 2382 46383 2614
rect 45809 2377 46383 2382
rect 13803 2075 13815 2307
rect 14021 2075 14032 2307
rect 13803 2059 14032 2075
rect 45808 2307 46384 2315
rect 45808 2075 45817 2307
rect 45903 2075 46289 2307
rect 46375 2075 46384 2307
rect 45808 2065 46384 2075
rect 53597 2307 53818 3112
rect 54492 2614 54854 3112
rect 54492 2382 54509 2614
rect 54836 2382 54854 2614
rect 54492 2361 54854 2382
rect 53597 2075 53614 2307
rect 53799 2075 53818 2307
rect 53597 2037 53818 2075
rect 164047 2307 164268 3112
rect 164942 2614 165304 3112
rect 164942 2382 164959 2614
rect 165286 2382 165304 2614
rect 164942 2361 165304 2382
rect 164047 2075 164064 2307
rect 164249 2075 164268 2307
rect 164047 2037 164268 2075
rect 227707 2307 227928 3113
rect 228602 2614 228964 3112
rect 228602 2382 228619 2614
rect 228946 2382 228964 2614
rect 228602 2361 228964 2382
rect 227707 2075 227724 2307
rect 227909 2075 227928 2307
rect 227707 2037 227928 2075
rect 232967 2307 233188 3112
rect 233862 2614 234220 3112
rect 233862 2382 233879 2614
rect 234206 2382 234220 2614
rect 233862 2361 234220 2382
rect 232967 2075 232984 2307
rect 233169 2075 233188 2307
rect 232967 2037 233188 2075
rect 236137 2307 236358 3112
rect 237032 2614 237390 3112
rect 237032 2382 237049 2614
rect 237376 2382 237390 2614
rect 237032 2361 237390 2382
rect 236137 2075 236154 2307
rect 236339 2075 236358 2307
rect 236137 2037 236358 2075
rect 238229 2307 238450 3112
rect 239124 2614 239482 3112
rect 239124 2382 239141 2614
rect 239468 2382 239482 2614
rect 239124 2361 239482 2382
rect 238229 2075 238246 2307
rect 238431 2075 238450 2307
rect 238229 2037 238450 2075
rect 240321 2307 240542 3112
rect 241216 2614 241574 3112
rect 241216 2382 241233 2614
rect 241560 2382 241574 2614
rect 241216 2361 241574 2382
rect 240321 2075 240338 2307
rect 240523 2075 240542 2307
rect 240321 2037 240542 2075
rect 242413 2307 242634 3112
rect 242768 2614 243126 3112
rect 242768 2382 242785 2614
rect 243112 2382 243126 2614
rect 242768 2361 243126 2382
rect 243197 2614 243436 3112
rect 243197 2382 243214 2614
rect 243386 2382 243436 2614
rect 243197 2361 243436 2382
rect 242413 2075 242430 2307
rect 242615 2075 242634 2307
rect 242413 2037 242634 2075
rect 243539 2307 243760 3112
rect 243881 2614 244124 3113
rect 243881 2382 243895 2614
rect 244112 2382 244124 2614
rect 243881 2362 244124 2382
rect 243539 2075 243556 2307
rect 243741 2075 243760 2307
rect 243539 2037 243760 2075
rect 244228 2307 244427 3114
rect 244228 2075 244239 2307
rect 244414 2075 244427 2307
rect 244228 2055 244427 2075
rect 12933 1912 13195 1940
rect 12933 1674 12943 1912
rect 13184 1674 13195 1912
rect 12933 -1873 13195 1674
rect 244859 1577 245137 1614
rect 244859 1343 244872 1577
rect 245127 1343 245137 1577
rect 45972 1236 46071 1304
rect 45972 677 45984 1236
rect 46053 677 46071 1236
rect 13297 -1526 45896 -1481
rect 13297 -1699 13322 -1526
rect 45823 -1699 45896 -1526
rect 13297 -1715 45896 -1699
rect 12933 -2111 12944 -1873
rect 13185 -1892 45896 -1873
rect 13185 -2065 13279 -1892
rect 45824 -2065 45896 -1892
rect 13185 -2111 45896 -2065
rect 12933 -4869 13195 -2111
rect 45972 -4207 46071 677
rect 244859 -1481 245137 1343
rect 46167 -1526 244871 -1481
rect 46167 -1700 46232 -1526
rect 244672 -1700 244871 -1526
rect 46167 -1715 244871 -1700
rect 245126 -1715 245137 -1481
rect 46167 -1889 244756 -1873
rect 46167 -2063 46232 -1889
rect 244672 -2063 244756 -1889
rect 46167 -2111 244756 -2063
rect 45972 -4774 45978 -4207
rect 46066 -4774 46071 -4207
rect 45972 -4780 46071 -4774
rect 12933 -5107 12944 -4869
rect 13185 -5107 13195 -4869
rect 244859 -5099 245137 -1715
rect 12933 -5141 13195 -5107
rect 12937 -5316 13077 -5308
rect 12937 -5504 12944 -5316
rect 13070 -5504 13077 -5316
rect 12937 -5776 13077 -5504
rect 23204 -5316 23425 -5278
rect 23204 -5504 23221 -5316
rect 23406 -5504 23425 -5316
rect 13534 -5572 13749 -5550
rect 13534 -5760 13541 -5572
rect 13741 -5760 13749 -5572
rect 13534 -5935 13749 -5760
rect 23204 -6353 23425 -5504
rect 69404 -5316 69625 -5278
rect 69404 -5504 69421 -5316
rect 69606 -5504 69625 -5316
rect 24099 -5572 24461 -5551
rect 24099 -5760 24116 -5572
rect 24443 -5760 24461 -5572
rect 24099 -6353 24461 -5760
rect 69404 -6353 69625 -5504
rect 122004 -5316 122225 -5277
rect 122004 -5504 122021 -5316
rect 122206 -5504 122225 -5316
rect 70299 -5572 70661 -5551
rect 70299 -5760 70316 -5572
rect 70643 -5760 70661 -5572
rect 70299 -6353 70661 -5760
rect 122004 -6352 122225 -5504
rect 174604 -5316 174825 -5277
rect 174604 -5504 174621 -5316
rect 174806 -5504 174825 -5316
rect 122899 -5572 123261 -5550
rect 122899 -5760 122916 -5572
rect 123243 -5760 123261 -5572
rect 122899 -6352 123261 -5760
rect 174604 -6352 174825 -5504
rect 227204 -5316 227425 -5277
rect 227204 -5504 227221 -5316
rect 227406 -5504 227425 -5316
rect 175499 -5572 175861 -5550
rect 175499 -5760 175516 -5572
rect 175843 -5760 175861 -5572
rect 175499 -6352 175861 -5760
rect 227204 -6352 227425 -5504
rect 244277 -5316 244411 -5300
rect 244277 -5504 244285 -5316
rect 244402 -5504 244411 -5316
rect 228099 -5572 228461 -5550
rect 228099 -5760 228116 -5572
rect 228443 -5760 228461 -5572
rect 228099 -6352 228461 -5760
rect 243887 -5572 244092 -5553
rect 243887 -5760 243897 -5572
rect 244079 -5760 244092 -5572
rect 243887 -6160 244092 -5760
rect 244277 -6158 244411 -5504
<< via3 >>
rect 13322 -1615 45823 -1526
rect 13322 -1699 45823 -1615
rect 13279 -1976 13323 -1892
rect 13323 -1976 45824 -1892
rect 13279 -2065 45824 -1976
rect 46232 -1615 244672 -1526
rect 46232 -1699 244671 -1615
rect 244671 -1699 244672 -1615
rect 46232 -1700 244672 -1699
rect 46232 -1890 244672 -1889
rect 46232 -1974 46233 -1890
rect 46233 -1974 244672 -1890
rect 46232 -2063 244672 -1974
<< metal4 >>
rect -892 -1526 245148 -33
rect -892 -1699 13322 -1526
rect 45823 -1699 46232 -1526
rect -892 -1700 46232 -1699
rect 244672 -1700 245148 -1526
rect -892 -1718 245148 -1700
rect -885 -1889 245155 -1869
rect -885 -1892 46232 -1889
rect -885 -2065 13279 -1892
rect 45824 -2063 46232 -1892
rect 244672 -2063 245155 -1889
rect 45824 -2065 245155 -2063
rect -885 -3554 245155 -2065
<< comment >>
rect 45874 -5615 45942 -5536
rect 46344 -5615 46412 -5536
rect 45874 -5773 46412 -5615
use bias_nstack  bias_nstack_0
array 0 439 -526 0 0 -3895
timestamp 1713991449
transform -1 0 17154 0 -1 -4733
box 3262 -2860 3922 1035
use bias_pstack  bias_pstack_0
array 0 439 526 0 0 -167
timestamp 1713995181
transform 1 0 11201 0 -1 -1327
box 1990 -3967 2710 388
use sky130_fd_pr__res_high_po_0p35_P35QVK  XR2 paramcells
timestamp 1713888873
transform 1 0 6139 0 1 -1753
box -6758 -3582 6758 3582
<< labels >>
flabel comment 46135 -5695 46135 -5695 0 FreeSans 1600 0 0 0 mirror
flabel metal2 46082 2684 46242 2884 0 FreeSans 256 0 0 0 enb
port 3 nsew
flabel metal3 227707 2872 227928 3113 0 FreeSans 1600 90 0 0 enb_600
port 17 nsew
flabel metal3 228602 2871 228964 3112 0 FreeSans 1600 90 0 0 src_600
port 18 nsew
flabel metal3 232967 2872 233188 3112 0 FreeSans 1600 90 0 0 enb_400
port 19 nsew
flabel metal3 233862 2872 234220 3112 0 FreeSans 1600 90 0 0 src_400
port 20 nsew
flabel metal3 236137 2872 236358 3112 0 FreeSans 1600 90 0 0 enb_200_0
port 21 nsew
flabel metal3 237032 2872 237390 3112 0 FreeSans 1600 90 0 0 src_200_0
port 22 nsew
flabel metal3 238229 2872 238450 3112 0 FreeSans 1600 90 0 0 enb_200_1
port 23 nsew
flabel metal3 239124 2872 239482 3112 0 FreeSans 1600 90 0 0 src_200_1
port 24 nsew
flabel metal3 240321 2872 240542 3112 0 FreeSans 1600 90 0 0 enb_200_2
port 25 nsew
flabel metal3 241216 2872 241574 3112 0 FreeSans 1600 90 0 0 src_200_2
port 26 nsew
flabel metal3 242413 2872 242634 3112 0 FreeSans 1600 90 0 0 enb_100
port 27 nsew
flabel metal3 242768 2872 243126 3112 0 FreeSans 1600 90 0 0 src_100
port 28 nsew
flabel metal3 53597 2897 53818 3112 0 FreeSans 1600 90 0 0 enb_10000_0
port 13 nsew
flabel metal3 54492 2871 54854 3112 0 FreeSans 1600 90 0 0 src_10000_0
port 14 nsew
flabel metal3 164047 2871 164268 3112 0 FreeSans 1600 90 0 0 enb_10000_1
port 16 nsew
flabel metal3 164942 2871 165304 3112 0 FreeSans 1600 90 0 0 src_10000_1
port 15 nsew
flabel metal3 69404 -6353 69625 -6124 0 FreeSans 1600 90 0 0 ena_5000_0
port 31 nsew
flabel metal3 122004 -6352 122225 -6123 0 FreeSans 1600 90 0 0 ena_5000_1
port 33 nsew
flabel metal3 174604 -6352 174825 -6123 0 FreeSans 1600 90 0 0 ena_5000_2
port 35 nsew
flabel metal1 -902 1231 -702 1431 0 FreeSans 256 0 0 0 ref_in
port 1 nsew
flabel metal3 243197 2872 243436 3112 0 FreeSans 1600 90 0 0 src_50
port 30 nsew
flabel metal3 243539 2872 243760 3112 0 FreeSans 1600 90 0 0 enb_50
port 29 nsew
flabel metal3 12937 -5776 13077 -5639 0 FreeSans 1600 90 0 0 ena_test0
port 39 nsew
flabel metal3 13534 -5935 13749 -5782 0 FreeSans 1600 90 0 0 snk_test0
port 40 nsew
flabel metal3 243887 -6160 244092 -6018 0 FreeSans 1600 90 0 0 snk_test1
port 41 nsew
flabel metal3 244277 -6158 244411 -6016 0 FreeSans 1600 90 0 0 ena_test1
port 42 nsew
flabel metal3 243881 2872 244124 3113 0 FreeSans 1600 90 0 0 src_test1
port 43 nsew
flabel metal3 244228 2873 244427 3114 0 FreeSans 1600 90 0 0 enb_test1
port 44 nsew
flabel metal3 13467 2695 13696 2928 0 FreeSans 1600 90 0 0 src_test0
port 45 nsew
flabel metal3 13803 2695 14032 2928 0 FreeSans 1600 90 0 0 enb_test0
port 46 nsew
flabel metal3 70299 -6353 70661 -6124 0 FreeSans 1600 90 0 0 snk_5000_0
port 48 nsew
flabel metal3 122899 -6352 123261 -6123 0 FreeSans 1600 90 0 0 snk_5000_1
port 34 nsew
flabel metal3 175499 -6352 175861 -6123 0 FreeSans 1600 90 0 0 snk_5000_2
port 36 nsew
flabel metal4 -892 -1718 -659 -33 0 FreeSans 1600 90 0 0 avdd
port 47 nsew
flabel metal4 -885 -3554 -652 -1869 0 FreeSans 1600 90 0 0 avss
port 12 nsew
flabel metal3 23204 -6353 23425 -6124 0 FreeSans 1600 90 0 0 ena_2000
port 49 nsew
flabel metal3 24099 -6353 24461 -6124 0 FreeSans 1600 90 0 0 snk_2000
port 32 nsew
flabel metal3 227204 -6352 227425 -6164 0 FreeSans 1600 90 0 0 ena_3700
port 38 nsew
flabel metal3 228099 -6352 228461 -6164 0 FreeSans 1600 90 0 0 snk_3700
port 37 nsew
flabel metal2 35144 -5790 35344 -5590 0 FreeSans 256 0 0 0 ena
port 11 nsew
<< end >>
