magic
tech sky130A
magscale 1 2
timestamp 1714090311
<< locali >>
rect 3392 364 3448 658
rect 3742 364 3926 658
rect 3392 342 3926 364
rect 3448 270 3742 342
<< metal1 >>
rect 3724 1027 3788 1035
rect 3568 771 3622 777
rect 3300 280 3352 290
rect 3352 144 3353 276
rect 3300 138 3353 144
rect 3301 -1916 3353 138
rect 3392 -1514 3456 52
rect 3568 -610 3622 583
rect 3724 -540 3788 839
rect 3834 282 3886 290
rect 3834 280 3887 282
rect 3886 144 3887 280
rect 3834 138 3887 144
rect 3568 -1622 3620 -860
rect 3301 -2632 3456 -1916
rect 3568 -2584 3620 -1818
rect 3726 -2502 3790 -936
rect 3568 -2586 3616 -2584
rect 3835 -2632 3887 138
rect 3301 -2690 3887 -2632
rect 3300 -2704 3890 -2690
rect 3300 -2782 3358 -2704
rect 3832 -2782 3890 -2704
rect 3300 -2796 3890 -2782
<< via1 >>
rect 3724 839 3788 1027
rect 3568 583 3622 771
rect 3300 144 3352 280
rect 3834 144 3886 280
rect 3568 -1818 3620 -1622
rect 3358 -2782 3832 -2704
<< metal2 >>
rect 3718 839 3724 1027
rect 3788 839 3794 1027
rect 3560 583 3568 771
rect 3622 583 3631 771
rect 3258 280 3926 374
rect 3258 144 3300 280
rect 3352 144 3834 280
rect 3886 144 3926 280
rect 3258 136 3926 144
rect 3258 -1622 3926 -1598
rect 3258 -1818 3568 -1622
rect 3620 -1818 3926 -1622
rect 3258 -1836 3926 -1818
rect 3258 -2704 3926 -2622
rect 3258 -2782 3358 -2704
rect 3832 -2782 3926 -2704
rect 3258 -2860 3926 -2782
use sky130_fd_pr__diode_pw2nd_05v5_FT76RK  sky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 paramcells
timestamp 1713888873
transform 1 0 3595 0 1 511
box -183 -183 183 183
use sky130_fd_pr__nfet_05v0_nvt_QRKT8P  XM6 paramcells
timestamp 1714090311
transform 1 0 3594 0 1 -1226
box -332 -558 332 558
use sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P  XM7 paramcells
timestamp 1714090311
transform 1 0 3594 0 1 -240
box -332 -558 332 558
use sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ  XM12 paramcells
timestamp 1714090311
transform 1 0 3594 0 1 -2212
box -332 -558 332 558
<< labels >>
flabel metal1 3724 690 3788 792 0 FreeSans 560 90 0 0 itail
port 2 nsew
flabel metal1 3568 404 3622 458 0 FreeSans 560 0 0 0 ena
port 3 nsew
flabel metal2 3262 -1836 3568 -1598 0 FreeSans 560 0 0 0 nbias
port 4 nsew
flabel metal1 3392 -612 3456 -550 0 FreeSans 560 90 0 0 vcasc
port 5 nsew
flabel metal2 3258 -2860 3358 -2622 0 FreeSans 560 90 0 0 avss
port 1 nsew
<< end >>
