magic
tech sky130A
timestamp 1714177271
<< pwell >>
rect -110 -110 110 110
<< mvpsubdiff >>
rect -92 86 92 92
rect -92 69 -38 86
rect 38 69 92 86
rect -92 63 92 69
rect -92 38 -63 63
rect -92 -38 -86 38
rect -69 -38 -63 38
rect 63 38 92 63
rect -92 -63 -63 -38
rect 63 -38 69 38
rect 86 -38 92 38
rect 63 -63 92 -38
rect -92 -69 92 -63
rect -92 -86 -38 -69
rect 38 -86 92 -69
rect -92 -92 92 -86
<< mvpsubdiffcont >>
rect -38 69 38 86
rect -86 -38 -69 38
rect 69 -38 86 38
rect -38 -86 38 -69
<< mvndiode >>
rect -24 18 24 24
rect -24 -18 -18 18
rect 18 -18 24 18
rect -24 -24 24 -18
<< mvndiodec >>
rect -18 -18 18 18
<< locali >>
rect -86 69 -38 86
rect 38 69 86 86
rect -86 38 -69 69
rect 69 38 86 69
rect -26 -18 -18 18
rect 18 -18 26 18
rect -86 -69 -69 -38
rect 69 -69 86 -38
rect -86 -86 -38 -69
rect 38 -86 86 -69
<< viali >>
rect -18 -18 18 18
<< metal1 >>
rect -24 18 24 21
rect -24 -18 -18 18
rect 18 -18 24 18
rect -24 -21 24 -18
<< properties >>
string FIXED_BBOX -77 -77 77 77
string gencell sky130_fd_pr__diode_pw2nd_11v0
string library sky130
string parameters w 0.48 l 0.48 area 230.399m peri 1.92 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
