* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_WHP78W a_131_6584# a_n367_6584# a_n1031_n7016#
+ a_961_n7016# a_n201_n7016# a_n699_n7016# a_n865_6584# a_463_n7016# a_463_6584# a_n699_6584#
+ a_n1197_6584# a_297_6584# a_1127_n7016# a_n533_n7016# a_961_6584# a_n35_n7016# a_795_n7016#
+ a_795_6584# a_n201_6584# a_629_6584# a_297_n7016# a_629_n7016# a_n35_6584# a_n865_n7016#
+ a_n1197_n7016# a_n367_n7016# a_n533_6584# a_n1327_n7146# a_131_n7016# a_n1031_6584#
+ a_1127_6584#
X0 a_n699_6584# a_n699_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X1 a_131_6584# a_131_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X2 a_n1197_6584# a_n1197_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X3 a_n533_6584# a_n533_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X4 a_1127_6584# a_1127_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X5 a_463_6584# a_463_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X6 a_629_6584# a_629_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X7 a_n1031_6584# a_n1031_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X8 a_n35_6584# a_n35_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X9 a_961_6584# a_961_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X10 a_n367_6584# a_n367_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X11 a_297_6584# a_297_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X12 a_n865_6584# a_n865_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X13 a_795_6584# a_795_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
X14 a_n201_6584# a_n201_n7016# a_n1327_n7146# sky130_fd_pr__res_xhigh_po_0p35 l=66
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_M35ED8 a_1210_n8616# a_546_8184# a_878_n8616#
+ a_n118_n8616# a_1210_8184# a_n450_8184# a_n1944_8184# a_n1778_n8616# a_1044_8184#
+ a_n284_8184# a_n948_n8616# a_n1778_8184# a_878_8184# a_380_n8616# a_1542_n8616#
+ a_712_n8616# a_2040_8184# a_n1280_n8616# a_2040_n8616# a_1542_8184# a_n118_8184#
+ a_n1612_n8616# a_n450_n8616# a_1044_n8616# a_214_n8616# a_n782_8184# a_1376_8184#
+ a_n1280_8184# a_n2110_n8616# a_380_8184# a_n1114_n8616# a_n616_8184# a_1874_n8616#
+ a_n1114_8184# a_48_n8616# a_214_8184# a_1874_8184# a_n1944_n8616# a_1376_n8616#
+ a_n782_n8616# a_546_n8616# a_n2110_8184# a_1708_n8616# a_1708_8184# a_48_8184# a_n1612_8184#
+ a_n1446_n8616# a_n2240_n8746# a_712_8184# a_n284_n8616# a_n948_8184# a_n616_n8616#
+ a_n1446_8184#
X0 a_n616_8184# a_n616_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X1 a_1044_8184# a_1044_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X2 a_546_8184# a_546_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X3 a_380_8184# a_380_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X4 a_n1114_8184# a_n1114_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X5 a_1708_8184# a_1708_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X6 a_1542_8184# a_1542_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X7 a_2040_8184# a_2040_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X8 a_n450_8184# a_n450_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X9 a_n1612_8184# a_n1612_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X10 a_n284_8184# a_n284_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X11 a_48_8184# a_48_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X12 a_n948_8184# a_n948_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X13 a_n782_8184# a_n782_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X14 a_1376_8184# a_1376_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X15 a_878_8184# a_878_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X16 a_n1446_8184# a_n1446_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X17 a_n2110_8184# a_n2110_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X18 a_1874_8184# a_1874_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X19 a_n1944_8184# a_n1944_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X20 a_214_8184# a_214_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X21 a_n1280_8184# a_n1280_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X22 a_1210_8184# a_1210_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X23 a_712_8184# a_712_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X24 a_n118_8184# a_n118_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
X25 a_n1778_8184# a_n1778_n8616# a_n2240_n8746# sky130_fd_pr__res_xhigh_po_0p35 l=82
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_VTNT3C a_n118_7484# a_214_n7916# a_48_n7916#
+ a_214_7484# a_n414_n8046# a_48_7484# a_n284_n7916# a_n118_n7916# a_n284_7484#
X0 a_n284_7484# a_n284_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
X1 a_48_7484# a_48_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
X2 a_214_7484# a_214_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
X3 a_n118_7484# a_n118_n7916# a_n414_n8046# sky130_fd_pr__res_xhigh_po_0p35 l=75
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_01v8_LHQHT5 a_n29_n400# a_887_n400# a_429_n400# a_n887_n488#
+ a_n1047_n574# a_n429_n488# a_487_n488# a_n945_n400# a_29_n488# a_n487_n400#
X0 a_n487_n400# a_n887_n488# a_n945_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X1 a_n29_n400# a_n429_n488# a_n487_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X2 a_429_n400# a_29_n488# a_n29_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X3 a_887_n400# a_487_n488# a_429_n400# a_n1047_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B a_29_n388# a_n129_n388# a_n321_n522# a_n29_n300#
+ a_n187_n300# a_129_n300#
X0 a_129_n300# a_29_n388# a_n29_n300# a_n321_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.5
X1 a_n29_n300# a_n129_n388# a_n187_n300# a_n321_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VHBZVD a_n400_n197# a_400_n100# w_n658_n397#
+ a_n458_n100#
X0 a_400_n100# a_n400_n197# a_n458_n100# w_n658_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt level_shift dvdd dvss in in_b out_b out dw_2668_n1758# avss avdd
XXM1 dvss in_b dvss in sky130_fd_pr__nfet_01v8_69TQ3K
XXM2 dvdd in dvdd in_b sky130_fd_pr__pfet_01v8_3HMWVM
XXM3 in in avss out_b avss avss sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
XXM4 in_b in_b avss out avss avss sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
XXM5 out avdd avdd out_b sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM6 out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
.ends

.subckt sky130_fd_pr__nfet_01v8_6G4XAN a_n29_n155# a_29_n243# a_n287_n155# a_n389_n329#
+ a_n229_n243# a_229_55# a_229_n155# a_n287_55# a_n29_55#
X0 a_n29_n155# a_n229_n243# a_n287_n155# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X1 a_229_n155# a_29_n243# a_n29_n155# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X2 a_229_55# a_29_n243# a_n29_55# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X3 a_n29_55# a_n229_n243# a_n287_55# a_n389_n329# sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
.ends

.subckt sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X17 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt ripple_dly_4 clkin ena doneb dvss dvdd
Xx1 clkin doneb dvss dvss dvdd dvdd x1/X sky130_fd_sc_hd__and2_0
Xx3 Qb1 Qb2 ena dvss dvss dvdd dvdd x3/Q Qb2 sky130_fd_sc_hd__dfrbp_1
Xx2 x1/X Qb1 ena dvss dvss dvdd dvdd x2/Q Qb1 sky130_fd_sc_hd__dfrbp_1
Xx4 Qb2 doneb ena dvss dvss dvdd dvdd x4/Q doneb sky130_fd_sc_hd__dfrbp_1
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
X0 VGND TE_B a_30_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Z A a_215_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0672 ps=0.85 w=0.64 l=0.15
X2 a_215_369# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.10855 ps=1.005 w=0.64 l=0.15
X3 a_215_47# a_30_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.07665 ps=0.785 w=0.42 l=0.15
X4 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR TE_B a_30_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.005 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_AHZR5K a_n458_n50# a_n400_n138# a_n560_n224# a_400_n50#
X0 a_400_n50# a_n400_n138# a_n458_n50# a_n560_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
.ends

.subckt ripl_dly_clk_buf clkin clkout ena stby stby_b dvdd dvss
Xx1 clkin ena ena_done_b dvss dvdd ripple_dly_4
Xx2 clkin stby_b stby_done_b dvss dvdd ripple_dly_4
Xx3 stby_b stby_done_b ena ena_done_b stby dvss dvss dvdd dvdd clk_disable sky130_fd_sc_hd__a221o_1
Xx5 clkin clk_disable dvss dvss dvdd dvdd clkout sky130_fd_sc_hd__einvn_0
XXM3 clkout clk_disable dvss dvss sky130_fd_pr__nfet_01v8_AHZR5K
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_68VL2P a_961_n11416# a_463_10984# a_n35_n11416#
+ a_1625_10984# a_n201_n11416# a_n1197_n11416# a_n1363_10984# a_1625_n11416# a_629_n11416#
+ a_1127_10984# a_131_n11416# a_n533_10984# a_n35_10984# a_n533_n11416# a_1957_n11416#
+ a_795_10984# a_n2157_n11546# a_463_n11416# a_1957_10984# a_n865_n11416# a_n1861_n11416#
+ a_n1695_10984# a_1791_n11416# a_1127_n11416# a_795_n11416# a_297_10984# a_1459_10984#
+ a_n865_10984# a_629_10984# a_n1529_n11416# a_n1031_n11416# a_n1197_10984# a_1459_n11416#
+ a_n1529_10984# a_n367_10984# a_n367_n11416# a_131_10984# a_n1363_n11416# a_n2027_10984#
+ a_297_n11416# a_1293_n11416# a_n699_n11416# a_n1031_10984# a_1791_10984# a_n1695_n11416#
+ a_961_10984# a_n201_10984# a_n2027_n11416# a_n699_10984# a_n1861_10984# a_1293_10984#
X0 a_1957_10984# a_1957_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X1 a_n1861_10984# a_n1861_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X2 a_463_10984# a_463_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X3 a_1791_10984# a_1791_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X4 a_n35_10984# a_n35_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X5 a_795_10984# a_795_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X6 a_n2027_10984# a_n2027_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X7 a_961_10984# a_961_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X8 a_n1197_10984# a_n1197_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X9 a_n1031_10984# a_n1031_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X10 a_1127_10984# a_1127_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X11 a_n1529_10984# a_n1529_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X12 a_n367_10984# a_n367_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X13 a_n201_10984# a_n201_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X14 a_1459_10984# a_1459_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X15 a_n1363_10984# a_n1363_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X16 a_n699_10984# a_n699_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X17 a_n533_10984# a_n533_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X18 a_1293_10984# a_1293_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X19 a_n1695_10984# a_n1695_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X20 a_297_10984# a_297_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X21 a_1625_10984# a_1625_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X22 a_n865_10984# a_n865_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X23 a_131_10984# a_131_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
X24 a_629_10984# a_629_n11416# a_n2157_n11546# sky130_fd_pr__res_xhigh_po_0p35 l=110
.ends

.subckt sky130_fd_pr__nfet_01v8_UY343Z a_n800_n138# a_n960_n224# a_n858_n50# a_800_n50#
X0 a_800_n50# a_n800_n138# a_n858_n50# a_n960_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_EDYT7U w_n996_n269# a_n858_n50# a_n800_n147# a_800_n50#
X0 a_800_n50# a_n800_n147# a_n858_n50# w_n996_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YG6WAD a_n287_n488# a_761_n400# a_819_n488# a_345_n488#
+ a_n1111_n622# a_n29_n400# a_n919_n488# a_n187_n400# a_n445_n488# a_503_n488# a_n819_n400#
+ a_n345_n400# a_n603_n488# a_661_n488# a_n977_n400# a_n761_n488# a_129_n400# a_n503_n400#
+ a_287_n400# a_n661_n400# a_919_n400# a_445_n400# a_29_n488# a_n129_n488# a_603_n400#
+ a_187_n488#
X0 a_n503_n400# a_n603_n488# a_n661_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n488# a_n187_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n488# a_445_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n819_n400# a_n919_n488# a_n977_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n661_n400# a_n761_n488# a_n819_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_919_n400# a_819_n488# a_761_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_n187_n400# a_n287_n488# a_n345_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_761_n400# a_661_n488# a_603_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_287_n400# a_187_n488# a_129_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_n345_n400# a_n445_n488# a_n503_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X10 a_129_n400# a_29_n488# a_n29_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X11 a_445_n400# a_345_n488# a_287_n400# a_n1111_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VMUSDZ m3_n2386_n11680# m3_n2386_2480# c1_n2346_n11640#
+ m3_n2386_n6960# m3_n2386_n2240# m3_n2386_7200#
X0 c1_n2346_n11640# m3_n2386_n11680# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X1 c1_n2346_n11640# m3_n2386_7200# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X2 c1_n2346_n11640# m3_n2386_n2240# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X3 c1_n2346_n11640# m3_n2386_2480# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
X4 c1_n2346_n11640# m3_n2386_n6960# sky130_fd_pr__cap_mim_m3_1 l=22 w=22
.ends

.subckt sky130_fd_pr__nfet_01v8_HZ6WG7 a_100_n75# a_n260_n249# a_n100_n163# a_n158_n75#
X0 a_100_n75# a_n100_n163# a_n158_n75# a_n260_n249# sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_67RTNB m3_n3798_n4520# c1_n3758_n4480#
X0 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X5 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X6 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X8 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X10 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 c1_n3758_n4480# m3_n3798_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WXTTNJ c1_n2146_n2000# m3_n2186_n2040#
X0 c1_n2146_n2000# m3_n2186_n2040# sky130_fd_pr__cap_mim_m3_1 l=20 w=20
.ends

.subckt sky130_fd_pr__diode_pd2nw_05v5_K4SERG a_n45_n45# w_n183_n183#
X0 a_n45_n45# w_n183_n183# sky130_fd_pr__diode_pd2nw_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GZN5JV a_208_n400# a_366_n400# a_n558_n622# a_108_n488#
+ a_50_n400# a_n208_n488# a_266_n488# a_n366_n488# a_n108_n400# a_n266_n400# a_n50_n488#
+ a_n424_n400#
X0 a_n266_n400# a_n366_n488# a_n424_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_366_n400# a_266_n488# a_208_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_50_n400# a_n50_n488# a_n108_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n108_n400# a_n208_n488# a_n266_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_208_n400# a_108_n488# a_50_n400# a_n558_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_F5PPB9 c1_n1946_n7680# m3_n1986_n3800# m3_n1986_4040#
+ m3_n1986_120# m3_n1986_n7720#
X0 c1_n1946_n7680# m3_n1986_n7720# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X1 c1_n1946_n7680# m3_n1986_120# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X2 c1_n1946_n7680# m3_n1986_4040# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X3 c1_n1946_n7680# m3_n1986_n3800# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E4RF2H a_2054_64# a_n2112_64# a_n1934_n961# a_898_n864#
+ a_n258_n864# a_778_n864# a_n1356_n961# a_898_64# a_n200_n961# a_n378_64# a_n956_64#
+ a_n1992_n864# a_2512_n864# a_2512_64# a_1534_n961# a_n2570_64# a_n1534_n864# a_2054_n864#
+ a_320_64# a_n1414_n864# a_956_n961# w_n2770_n1161# a_n778_n961# a_1476_64# a_778_64#
+ a_n1534_64# a_n2512_n961# a_n258_64# a_n836_64# a_378_n961# a_320_n864# a_n956_n864#
+ a_1934_n864# a_200_64# a_200_n864# a_n2570_n864# a_1476_n864# a_n836_n864# a_1934_64#
+ a_1356_64# a_n1414_64# a_2112_n961# a_n378_n864# a_n1992_64# a_1356_n864# a_n2112_n864#
X0 a_n2112_64# a_n2512_n961# a_n2570_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X1 a_n2112_n864# a_n2512_n961# a_n2570_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X2 a_n1534_n864# a_n1934_n961# a_n1992_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X3 a_200_n864# a_n200_n961# a_n258_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X4 a_1356_n864# a_956_n961# a_898_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X5 a_778_64# a_378_n961# a_320_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X6 a_n956_64# a_n1356_n961# a_n1414_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X7 a_n956_n864# a_n1356_n961# a_n1414_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X8 a_1356_64# a_956_n961# a_898_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X9 a_1934_64# a_1534_n961# a_1476_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X10 a_778_n864# a_378_n961# a_320_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X11 a_n1534_64# a_n1934_n961# a_n1992_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X12 a_200_64# a_n200_n961# a_n258_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X13 a_n378_n864# a_n778_n961# a_n836_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X14 a_2512_n864# a_2112_n961# a_2054_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X15 a_n378_64# a_n778_n961# a_n836_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X16 a_1934_n864# a_1534_n961# a_1476_n864# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X17 a_2512_64# a_2112_n961# a_2054_64# w_n2770_n1161# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_74GBJT a_n208_n497# a_266_n497# a_208_n400# a_n366_n497#
+ a_366_n400# a_n50_n497# a_50_n400# a_n108_n400# a_n266_n400# w_n624_n697# a_n424_n400#
+ a_108_n497#
X0 a_n266_n400# a_n366_n497# a_n424_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_366_n400# a_266_n497# a_208_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_50_n400# a_n50_n497# a_n108_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n108_n400# a_n208_n497# a_n266_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_208_n400# a_108_n497# a_50_n400# w_n624_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_3H68VM w_n296_n619# a_n100_n497# a_100_n400# a_n158_n400#
X0 a_100_n400# a_n100_n497# a_n158_n400# w_n296_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6RLJVT a_n50_n497# a_50_n400# w_n308_n697# a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_MTZJAC a_761_n400# a_n29_n400# a_n187_n400# a_n819_n400#
+ a_n345_n400# a_29_n497# a_n129_n497# a_187_n497# a_129_n400# a_n503_n400# a_n287_n497#
+ a_287_n400# a_n661_n400# a_345_n497# a_n445_n497# a_445_n400# a_503_n497# a_n603_n497#
+ a_661_n497# w_n957_n619# a_603_n400# a_n761_n497#
X0 a_n661_n400# a_n761_n497# a_n819_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_n187_n400# a_n287_n497# a_n345_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_761_n400# a_661_n497# a_603_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X3 a_287_n400# a_187_n497# a_129_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_n345_n400# a_n445_n497# a_n503_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_129_n400# a_29_n497# a_n29_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X6 a_445_n400# a_345_n497# a_287_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n503_n400# a_n603_n497# a_n661_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_n29_n400# a_n129_n497# a_n187_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_603_n400# a_503_n497# a_445_n400# w_n957_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_Z6W9J4 a_2223_n200# a_n1703_n200# a_1245_n288#
+ a_n1245_n200# a_n1125_n200# a_667_n288# a_n489_n288# a_n2223_n288# a_1765_n200#
+ a_n667_n200# a_89_n288# a_1645_n200# a_31_n200# a_n2281_n200# a_1187_n200# a_n547_n200#
+ a_1067_n200# a_n89_n200# a_n1645_n288# a_609_n200# a_489_n200# a_1823_n288# a_n1067_n288#
+ a_n1823_n200# a_n2415_n422#
X0 a_n89_n200# a_n489_n288# a_n547_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X1 a_1645_n200# a_1245_n288# a_1187_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X2 a_n1823_n200# a_n2223_n288# a_n2281_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X3 a_n1245_n200# a_n1645_n288# a_n1703_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X4 a_489_n200# a_89_n288# a_31_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X5 a_1067_n200# a_667_n288# a_609_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X6 a_n667_n200# a_n1067_n288# a_n1125_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X7 a_2223_n200# a_1823_n288# a_1765_n200# a_n2415_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8CDM6Z a_n887_n497# a_n29_n400# w_n1145_n697#
+ a_887_n400# a_n429_n497# a_487_n497# a_429_n400# a_29_n497# a_n945_n400# a_n487_n400#
X0 a_n487_n400# a_n887_n497# a_n945_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X1 a_n29_n400# a_n429_n497# a_n487_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X2 a_429_n400# a_29_n497# a_n29_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=2
X3 a_887_n400# a_487_n497# a_429_n400# w_n1145_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_UYSCL3 c1_n1852_n1560# m3_n1892_120# m3_n150_130#
+ c1_n110_n1550# m3_n150_n1590# m3_n1892_n1600#
X0 c1_n110_n1550# m3_n150_n1590# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1 c1_n1852_n1560# m3_n1892_120# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X2 c1_n1852_n1560# m3_n1892_n1600# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X3 c1_n110_n1550# m3_n150_130# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_43FTN9 m3_n3546_n7996# c1_n3506_n7956#
X0 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X5 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X6 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X8 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X10 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X12 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X13 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X14 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X15 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X16 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X17 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X18 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X20 c1_n3506_n7956# m3_n3546_n7996# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_3DMTNZ m3_n2492_120# m3_n134_n2252# m3_n136_122#
+ c1_n2452_160# m3_n2490_n2254#
X0 c1_n2452_160# m3_n2492_120# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n2452_160# m3_n2490_n2254# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n2452_160# m3_n134_n2252# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n2452_160# m3_n136_122# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4HHTN9 m3_n1186_n4520# c1_n1146_n4480#
X0 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__pfet_01v8_M6QFHF a_229_n164# a_229_64# a_n287_64# a_n29_64#
+ a_29_n261# a_n29_n164# a_n229_n261# w_n425_n383# a_n287_n164#
X0 a_n29_64# a_n229_n261# a_n287_64# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X1 a_n29_n164# a_n229_n261# a_n287_n164# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=1
X2 a_229_n164# a_29_n261# a_n29_n164# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
X3 a_229_64# a_29_n261# a_n29_64# w_n425_n383# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H6M2KM a_n2516_n42# a_2458_n42# a_800_n42# a_858_n130#
+ a_n2650_n264# a_n800_n130# a_n2458_n130#
X0 a_800_n42# a_n800_n130# a_n858_n42# a_n2650_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X1 a_n858_n42# a_n2458_n130# a_n2516_n42# a_n2650_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X2 a_2458_n42# a_858_n130# a_800_n42# a_n2650_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_BKL7UB a_n1414_n855# a_n1548_n1077# a_778_55#
+ a_n836_55# a_n258_55# a_n1356_n943# a_n200_n943# a_320_n855# a_n956_n855# a_200_55#
+ a_200_n855# a_n836_n855# a_n1414_55# a_1356_55# a_n378_n855# a_1356_n855# a_956_n943#
+ a_n778_n943# a_898_n855# a_n258_n855# a_778_n855# a_378_n943# a_898_55# a_n956_55#
+ a_n378_55# a_320_55#
X0 a_n956_55# a_n1356_n943# a_n1414_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X1 a_n956_n855# a_n1356_n943# a_n1414_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X2 a_1356_55# a_956_n943# a_898_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X3 a_778_n855# a_378_n943# a_320_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X4 a_200_55# a_n200_n943# a_n258_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X5 a_n378_n855# a_n778_n943# a_n836_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X6 a_n378_55# a_n778_n943# a_n836_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X7 a_200_n855# a_n200_n943# a_n258_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X8 a_1356_n855# a_956_n943# a_898_n855# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
X9 a_778_55# a_378_n943# a_320_55# a_n1548_n1077# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_Y7GPAW a_n287_n488# a_761_n400# a_345_n488# a_n29_n400#
+ a_n187_n400# a_n445_n488# a_503_n488# a_n819_n400# a_n345_n400# a_n603_n488# a_661_n488#
+ a_n761_n488# a_129_n400# a_n503_n400# a_287_n400# a_n661_n400# a_n921_n574# a_445_n400#
+ a_29_n488# a_n129_n488# a_603_n400# a_187_n488#
X0 a_n503_n400# a_n603_n488# a_n661_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n488# a_n187_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n488# a_445_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n661_n400# a_n761_n488# a_n819_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n187_n400# a_n287_n488# a_n345_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_761_n400# a_661_n488# a_603_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_287_n400# a_187_n488# a_129_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n345_n400# a_n445_n488# a_n503_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_129_n400# a_29_n488# a_n29_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_445_n400# a_345_n488# a_287_n400# a_n921_n574# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_LL48TN a_n1802_n464# a_86_n561# a_2202_n464# a_1744_64#
+ a_n1802_64# a_486_64# a_n544_n464# a_n1116_n464# a_n544_64# a_658_n561# a_600_n464#
+ a_1172_64# a_n86_64# a_n1230_64# a_1630_n464# a_n1688_n464# a_28_64# a_1172_n464#
+ a_n86_n464# a_n2202_n561# a_n1688_64# a_1058_64# a_n1116_64# a_n658_n464# a_1744_n464#
+ a_486_n464# a_n1630_n561# w_n2398_n683# a_1630_64# a_1058_n464# a_n2260_n464# a_28_n464#
+ a_n658_64# a_1230_n561# a_n1230_n464# a_n1058_n561# a_n486_n561# a_600_64# a_2202_64#
+ a_1802_n561# a_n2260_64#
X0 a_1058_64# a_658_n561# a_600_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X1 a_2202_64# a_1802_n561# a_1744_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X2 a_n1802_n464# a_n2202_n561# a_n2260_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X3 a_486_n464# a_86_n561# a_28_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X4 a_1630_64# a_1230_n561# a_1172_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X5 a_486_64# a_86_n561# a_28_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X6 a_n1802_64# a_n2202_n561# a_n2260_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X7 a_1058_n464# a_658_n561# a_600_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X8 a_2202_n464# a_1802_n561# a_1744_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X9 a_n1230_n464# a_n1630_n561# a_n1688_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X10 a_1630_n464# a_1230_n561# a_1172_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X11 a_n86_64# a_n486_n561# a_n544_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X12 a_n658_n464# a_n1058_n561# a_n1116_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X13 a_n86_n464# a_n486_n561# a_n544_n464# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X14 a_n1230_64# a_n1630_n561# a_n1688_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
X15 a_n658_64# a_n1058_n561# a_n1116_64# w_n2398_n683# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_be_ip__lsxo avdd dvdd ibias ena standby dout xout xin avss_ip dvss_ip
+ avss dvss
Xamp_XR1 m1_24220_n8834# m1_24220_n8502# m1_10618_n7674# m1_10620_n9664# m1_10620_n8670#
+ m1_10620_n8006# m1_24220_n7840# m1_10620_n9334# m1_24220_n9166# m1_24220_n8172#
+ inv_in m1_24220_n9166# li_9150_n9268# m1_10620_n8338# m1_24220_n9832# m1_10620_n8670#
+ m1_10620_n9664# m1_24220_n9500# m1_24220_n8502# m1_24220_n9500# m1_10620_n9002#
+ m1_10620_n9334# m1_24220_n8834# m1_10620_n8006# m1_10618_n7674# m1_10620_n8338#
+ m1_24220_n8172# dvss_ip m1_10620_n9002# m1_24220_n7840# m1_24220_n9832# sky130_fd_pr__res_xhigh_po_0p35_WHP78W
Xbias_XR2 m1_2130_n17240# m1_18932_n16742# m1_2130_n16908# m1_2132_n15912# m1_18932_n17406#
+ m1_18932_n15746# vg2 m1_2132_n14254# m1_18932_n17074# m1_18932_n15746# m1_2132_n15248#
+ m1_18932_n14418# m1_18932_n17074# m1_2132_n16576# m1_2132_n17570# m1_2130_n16908#
+ avss_ip m1_2132_n14916# avss_ip m1_18932_n17738# m1_18932_n16078# m1_2134_n14584#
+ m1_2130_n15578# m1_2130_n17240# m1_2132_n16242# m1_18932_n15414# m1_18932_n17406#
+ m1_18932_n14750# avss_ip m1_18932_n16410# m1_2132_n14916# m1_18932_n15414# m1_2132_n17904#
+ m1_18932_n15082# m1_2132_n16242# m1_18932_n16410# vg1 m1_2132_n14254# m1_2132_n17570#
+ m1_2132_n15248# m1_2132_n16576# avss_ip m1_2132_n17904# m1_18932_n17738# m1_18932_n16078#
+ m1_18932_n14418# m1_2134_n14584# avss_ip m1_18932_n16742# m1_2132_n15912# m1_18932_n15082#
+ m1_2130_n15578# m1_18932_n14750# sky130_fd_pr__res_xhigh_po_0p35_M35ED8
Xx1 ena dvss dvss dvdd dvdd ena_ip sky130_fd_sc_hd__buf_1
Xbias_XR3 avss_ip avss_ip m1_3134_n13314# avss_ip avss_ip vrb avss_ip m1_3134_n13314#
+ avss_ip sky130_fd_pr__res_xhigh_po_0p35_VTNT3C
Xesd_n_xout avss_ip xout sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xx2 standby dvss dvss dvdd dvdd standby_ip sky130_fd_sc_hd__buf_1
Xant_diode_standby dvss standby sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xamp_XM4_18 dvss_ip xin_buf xin_buf vn dvss_ip vn vn vn vn vn sky130_fd_pr__nfet_01v8_LHQHT5
Xx3 dvdd dvss ena_ip x3/in_b x3/out_b x3/out avdd avss avdd level_shift
Xx4 dvdd dvss standby_ip standby_b x4/out_b standby_33 avdd avss avdd level_shift
Xesd_n_xin avss_ip xin sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xamp_XM11_13 dvss_ip inv_m2 inv_m2 dvss_ip inv_m1 dout_ip dout_ip dvss_ip dvss_ip
+ sky130_fd_pr__nfet_01v8_6G4XAN
Xx7 dout_ip dout_filt ena_ip standby_ip standby_b dvdd dvss ripl_dly_clk_buf
Xbias_XM5 icnode avss_ip avss_ip vg2 sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXR2 m1_2130_n21506# m1_24530_n21008# m1_2130_n20510# m1_24528_n22338# m1_2130_n20510#
+ m1_2130_n19514# m1_24530_n19348# m1_2128_n22170# m1_2128_n21174# m1_24530_n21672#
+ m1_2130_n20842# m1_24530_n20012# m1_24530_n20676# m1_2130_n20180# avss_ip m1_24528_n21342#
+ avss_ip m1_2128_n21174# avss_ip m1_2130_n19846# m1_2130_n18850# m1_24530_n19016#
+ xin m1_2130_n21838# m1_2130_n21506# m1_24530_n21008# m1_24528_n22004# m1_24530_n19680#
+ m1_24528_n21342# m1_2130_n19184# m1_2130_n19514# m1_24530_n19348# m1_2128_n22170#
+ m1_24530_n19016# m1_24530_n20344# m1_2130_n20180# m1_24530_n20676# m1_2130_n19184#
+ avss_ip m1_2130_n20842# m1_2130_n21838# m1_2130_n19846# m1_24530_n19680# m1_24528_n22338#
+ m1_2130_n18850# m1_24530_n21672# m1_24530_n20344# avss_ip m1_24530_n20012# xout
+ m1_24528_n22004# sky130_fd_pr__res_xhigh_po_0p35_68VL2P
Xamp_XM7 inv_in dvss_ip inv_m1 dvss_ip sky130_fd_pr__nfet_01v8_UY343Z
Xamp_XM6 dvdd_ip inv_m1 inv_in dvdd_ip sky130_fd_pr__pfet_01v8_EDYT7U
Xamp_XM8 dvdd_ip dvdd_ip li_9150_n9268# li_9150_n9268# sky130_fd_pr__pfet_01v8_EDYT7U
XXM1 xin avss_ip xin xin avss_ip xout xin avss_ip xin xin avss_ip xout xin xin avss_ip
+ xin avss_ip avss_ip xout xout avss_ip avss_ip xin xin xout xin sky130_fd_pr__nfet_g5v0d10v5_YG6WAD
Xamp_XM9 li_9150_n9268# dvss_ip li_9150_n9268# dvss_ip sky130_fd_pr__nfet_01v8_UY343Z
XXM3 dvss standby_ip dvss dout_ip sky130_fd_pr__nfet_01v8_AHZR5K
Xbias_XC1 xin xin vg1 xin xin xin sky130_fd_pr__cap_mim_m3_1_VMUSDZ
XXM4 dout dvss_ip dout_filt dvss_ip sky130_fd_pr__nfet_01v8_HZ6WG7
Xamp_XC1 xin_buf inv_in sky130_fd_pr__cap_mim_m3_1_67RTNB
Xbias_XC2 avdd_ip icnode sky130_fd_pr__cap_mim_m3_1_WXTTNJ
Xesd_p_xout xout avdd_ip sky130_fd_pr__diode_pd2nw_05v5_K4SERG
XXM5 avss_ip avss avss x3/out avss x3/out x3/out x3/out avss_ip avss x3/out avss_ip
+ sky130_fd_pr__nfet_g5v0d10v5_GZN5JV
Xbias_XC3 avss_ip vg2 vg2 vg2 vg2 sky130_fd_pr__cap_mim_m3_1_F5PPB9
XXM2_bias_XM3_4 avdd_ip avdd_ip vbreg avdd_ip li_22598_n15512# avdd_ip vbreg avdd_ip
+ vbreg xout avdd_ip avdd_ip avdd_ip avdd_ip vbreg avdd_ip xout avdd_ip xout xout
+ vbreg avdd_ip vbreg xout avdd_ip xout vbreg xout avdd_ip vbreg vbreg avdd_ip avdd_ip
+ xout li_22598_n15512# avdd_ip xout avdd_ip avdd_ip xout xout vbreg vg1 avdd_ip xout
+ avdd_ip sky130_fd_pr__pfet_g5v0d10v5_E4RF2H
Xant_diode_ena dvss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXM6 x3/out_b x3/out_b avdd_ip x3/out_b avdd x3/out_b avdd avdd_ip avdd avdd avdd_ip
+ x3/out_b sky130_fd_pr__pfet_g5v0d10v5_74GBJT
XXM7 dvdd_ip dout_filt dout dvdd_ip sky130_fd_pr__pfet_01v8_3H68VM
XXM9 standby_33 ibias ibias ibias_ip sky130_fd_pr__pfet_g5v0d10v5_6RLJVT
XXM8 dvdd dvdd_ip dvdd dvdd dvdd_ip standby_ip standby_ip standby_ip dvdd dvdd standby_ip
+ dvdd_ip dvdd_ip standby_ip standby_ip dvdd standby_ip standby_ip standby_ip dvdd
+ dvdd_ip standby_ip sky130_fd_pr__pfet_01v8_MTZJAC
Xamp_XM1_2 dvss_ip dvss_ip ibias_ip ibias_ip ibias_ip ibias_ip ibias_ip ibias_ip dvss_ip
+ dvss_ip ibias_ip dvss_ip vbp dvss_ip ibias_ip dvss_ip ibias_ip ibias_ip ibias_ip
+ dvss_ip dvss_ip ibias_ip ibias_ip dvss_ip dvss_ip sky130_fd_pr__nfet_g5v0d10v5_Z6W9J4
Xamp_XM3_5 xin tail dvdd_ip xin_buf xin xout xin_buf xout vn vn sky130_fd_pr__pfet_g5v0d10v5_8CDM6Z
Xesd_p_xin xin avdd_ip sky130_fd_pr__diode_pd2nw_05v5_K4SERG
XXC1 avdd_ip avss_ip avss_ip avdd_ip avss_ip avss_ip sky130_fd_pr__cap_mim_m3_1_UYSCL3
XXC2 dvss_ip dvdd_ip sky130_fd_pr__cap_mim_m3_1_43FTN9
XXC3 avdd avdd avdd avss avdd sky130_fd_pr__cap_mim_m3_1_3DMTNZ
XXC4 dvss dvdd sky130_fd_pr__cap_mim_m3_1_4HHTN9
Xamp_XM10_12 dout_ip dout_ip inv_m2 dvdd_ip inv_m2 dvdd_ip inv_m1 dvdd_ip dvdd_ip
+ sky130_fd_pr__pfet_01v8_M6QFHF
Xbias_XM6_7_8 vbreg avss_ip li_8336_n12442# li_8336_n12442# avss_ip icnode icnode
+ sky130_fd_pr__nfet_g5v0d10v5_H6M2KM
Xbias_XM1_2 avss_ip avss_ip vrb vrb avss_ip avss_ip vg1 vbreg avss_ip vg1 vbreg vrb
+ avss_ip avss_ip vbreg avss_ip avss_ip vg2 avss_ip vbreg vrb vg2 avss_ip avss_ip
+ vbreg vbreg sky130_fd_pr__nfet_g5v0d10v5_BKL7UB
XXM11 standby_b dvss standby_b dvss_ip dvss standby_b standby_b dvss dvss_ip standby_b
+ standby_b standby_b dvss dvss dvss_ip dvss_ip dvss dvss standby_b standby_b dvss_ip
+ standby_b sky130_fd_pr__nfet_01v8_Y7GPAW
Xamp_XM16_17 dvdd_ip vbp dvdd_ip dvdd_ip dvdd_ip dvdd_ip dvdd_ip tail dvdd_ip vbp
+ dvdd_ip tail dvdd_ip tail dvdd_ip dvdd_ip vbp tail tail vbp dvdd_ip tail tail dvdd_ip
+ dvdd_ip dvdd_ip vbp dvdd_ip dvdd_ip tail dvdd_ip tail dvdd_ip vbp tail vbp vbp dvdd_ip
+ dvdd_ip vbp dvdd_ip sky130_fd_pr__pfet_01v8_LL48TN
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RK a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_QRKT8P a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_05v0_nvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_nstack itail ena nbias avss vcasc
XXM12 avss avss nbias m1_3726_n2502# sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RK
XXM6 avss vcasc nbias m1_3726_n2502# sky130_fd_pr__nfet_05v0_nvt_QRKT8P
XXM7 avss vcasc ena itail sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P
.ends

.subckt sky130_fd_pr__res_high_po_0p35_P35QVK a_380_2984# a_5692_n3416# a_n3770_2984#
+ a_3866_2984# a_3202_n3416# a_n1446_n3416# a_n284_n3416# a_n616_2984# a_4696_n3416#
+ a_4198_2984# a_2206_n3416# a_n1114_2984# a_n4102_2984# a_n616_n3416# a_6190_n3416#
+ a_n6592_2984# a_2372_2984# a_n5762_n3416# a_5360_2984# a_214_2984# a_n3604_2984#
+ a_1210_n3416# a_5194_n3416# a_6522_n3416# a_n4766_n3416# a_1874_2984# a_4862_2984#
+ a_4198_n3416# a_5526_n3416# a_5194_2984# a_n6260_n3416# a_878_n3416# a_n3438_2984#
+ a_n2110_2984# a_n6426_2984# a_2206_2984# a_n118_n3416# a_n3770_n3416# a_4696_2984#
+ a_n5264_n3416# a_48_2984# a_4530_n3416# a_n2774_n3416# a_n1612_2984# a_n4600_2984#
+ a_n5928_2984# a_1708_2984# a_6024_n3416# a_n4268_n3416# a_2870_2984# a_3534_n3416#
+ a_712_2984# a_n1778_n3416# a_5028_2984# a_5028_n3416# a_n948_2984# a_2538_n3416#
+ a_6190_2984# a_n1446_2984# a_n3272_n3416# a_n4434_2984# a_n4600_n3416# a_3202_2984#
+ a_n948_n3416# a_5692_2984# a_380_n3416# a_546_2984# a_4032_n3416# a_n2276_n3416#
+ a_n3604_n3416# a_n3936_2984# a_1542_n3416# a_2704_2984# a_3036_n3416# a_712_n3416#
+ a_n2608_n3416# a_n4268_2984# a_3036_2984# a_6024_2984# a_5858_n3416# a_n1280_n3416#
+ a_n6592_n3416# a_n2442_2984# a_n4102_n3416# a_2538_2984# a_n5430_2984# a_2040_n3416#
+ a_5526_2984# a_1210_2984# a_n1612_n3416# a_n5596_n3416# a_4862_n3416# a_n450_n3416#
+ a_n1944_2984# a_n3106_n3416# a_n4932_2984# a_1044_n3416# a_n450_2984# a_3700_2984#
+ a_6356_n3416# a_214_n3416# a_n5928_n3416# a_n6722_n3546# a_3866_n3416# a_n2276_2984#
+ a_n5264_2984# a_1044_2984# a_4032_2984# a_n2110_n3416# a_n6094_n3416# a_n1778_2984#
+ a_n4766_2984# a_5360_n3416# a_n284_2984# a_3534_2984# a_n4932_n3416# a_6522_2984#
+ a_n1114_n3416# a_2870_n3416# a_n5098_n3416# a_n6426_n3416# a_878_2984# a_4364_n3416#
+ a_n5098_2984# a_n3936_n3416# a_n2940_2984# a_1874_n3416# a_3368_n3416# a_n3272_2984#
+ a_3368_2984# a_48_n3416# a_n6260_2984# a_2040_2984# a_6356_2984# a_n5430_n3416#
+ a_n2940_n3416# a_n118_2984# a_n2774_2984# a_n4434_n3416# a_n5762_2984# a_1542_2984#
+ a_2372_n3416# a_4530_2984# a_5858_2984# a_3700_n3416# a_n1944_n3416# a_n3438_n3416#
+ a_n6094_2984# a_n782_n3416# a_1376_n3416# a_n782_2984# a_2704_n3416# a_546_n3416#
+ a_n3106_2984# a_n1280_2984# a_n5596_2984# a_1376_2984# a_1708_n3416# a_4364_2984#
+ a_n2442_n3416# a_n2608_2984#
X0 a_n3936_2984# a_n3936_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X1 a_n1612_2984# a_n1612_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X2 a_n6592_2984# a_n6592_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X3 a_n4434_2984# a_n4434_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X4 a_48_2984# a_48_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X5 a_2704_2984# a_2704_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X6 a_4862_2984# a_4862_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X7 a_3202_2984# a_3202_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X8 a_5360_2984# a_5360_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X9 a_5526_2984# a_5526_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X10 a_n948_2984# a_n948_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X11 a_n782_2984# a_n782_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X12 a_6024_2984# a_6024_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X13 a_n4932_2984# a_n4932_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X14 a_1376_2984# a_1376_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X15 a_878_2984# a_878_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X16 a_4198_2984# a_4198_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X17 a_n3770_2984# a_n3770_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X18 a_n1446_2984# a_n1446_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X19 a_3700_2984# a_3700_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X20 a_n4268_2984# a_n4268_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X21 a_n2110_2984# a_n2110_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X22 a_1874_2984# a_1874_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X23 a_6522_2984# a_6522_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X24 a_2372_2984# a_2372_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X25 a_2538_2984# a_2538_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X26 a_4696_2984# a_4696_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X27 a_3036_2984# a_3036_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X28 a_5194_2984# a_5194_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X29 a_n1944_2984# a_n1944_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X30 a_n4766_2984# a_n4766_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X31 a_n2608_2984# a_n2608_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X32 a_n2442_2984# a_n2442_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X33 a_214_2984# a_214_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X34 a_n5430_2984# a_n5430_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X35 a_n5264_2984# a_n5264_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X36 a_n3106_2984# a_n3106_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X37 a_2870_2984# a_2870_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X38 a_n1280_2984# a_n1280_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X39 a_1210_2984# a_1210_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X40 a_3534_2984# a_3534_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X41 a_5692_2984# a_5692_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X42 a_5858_2984# a_5858_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X43 a_712_2984# a_712_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X44 a_4032_2984# a_4032_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X45 a_6190_2984# a_6190_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X46 a_6356_2984# a_6356_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X47 a_n5928_2984# a_n5928_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X48 a_n5762_2984# a_n5762_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X49 a_n3604_2984# a_n3604_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X50 a_n118_2984# a_n118_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X51 a_n6426_2984# a_n6426_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X52 a_n4102_2984# a_n4102_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X53 a_n1778_2984# a_n1778_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X54 a_4530_2984# a_4530_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X55 a_n4600_2984# a_n4600_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X56 a_n2276_2984# a_n2276_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X57 a_n5098_2984# a_n5098_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X58 a_n616_2984# a_n616_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X59 a_1044_2984# a_1044_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X60 a_3368_2984# a_3368_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X61 a_546_2984# a_546_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X62 a_n2940_2984# a_n2940_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X63 a_n2774_2984# a_n2774_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X64 a_380_2984# a_380_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X65 a_n5596_2984# a_n5596_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X66 a_n3438_2984# a_n3438_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X67 a_n3272_2984# a_n3272_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X68 a_n1114_2984# a_n1114_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X69 a_n6260_2984# a_n6260_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X70 a_n6094_2984# a_n6094_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X71 a_1708_2984# a_1708_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X72 a_1542_2984# a_1542_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X73 a_2206_2984# a_2206_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X74 a_3866_2984# a_3866_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X75 a_2040_2984# a_2040_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X76 a_4364_2984# a_4364_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X77 a_5028_2984# a_5028_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X78 a_n450_2984# a_n450_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X79 a_n284_2984# a_n284_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ a_n158_n300# w_n362_n597# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n362_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_H75TTW a_n158_n300# w_n362_n597# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n362_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_pstack pcasc enb itail vcasc pbias avss avdd
XXM13 m1_2150_n1558# avdd pcasc vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__pfet_g5v0d10v5_G8LMTZ_0 itail avdd enb vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss enb sky130_fd_pr__diode_pw2nd_05v5_FT76RK
Xsky130_fd_pr__pfet_g5v0d10v5_H75TTW_0 m1_2150_n1558# avdd pbias avdd sky130_fd_pr__pfet_g5v0d10v5_H75TTW
.ends

.subckt bias_generator ref_in enb ena enb_10000_0 src_10000_0 src_10000_1 enb_10000_1
+ enb_600 src_600 enb_400 src_400 enb_200_0 src_200_0 enb_200_1 src_200_1 enb_200_2
+ src_200_2 enb_100 src_100 enb_50 src_50 ena_5000_0 snk_2000 snk_5000_1 ena_5000_2
+ snk_5000_2 snk_3700 ena_3700 ena_test0 snk_test0 snk_test1 ena_test1 src_test1 enb_test1
+ src_test0 enb_test0 snk_5000_0 ena_2000 vsub ena_5000_1 avdd avss
Xbias_nstack_0[0] snk_test0 ena_test0 bias_nstack_0[9]/nbias avss bias_nstack_0[0]/vcasc
+ bias_nstack
Xbias_nstack_0[1] snk_test0 ena_test0 bias_nstack_0[9]/nbias avss bias_nstack_0[1]/vcasc
+ bias_nstack
Xbias_nstack_0[2] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[2]/vcasc
+ bias_nstack
Xbias_nstack_0[3] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[3]/vcasc
+ bias_nstack
Xbias_nstack_0[4] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[4]/vcasc
+ bias_nstack
Xbias_nstack_0[5] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[5]/vcasc
+ bias_nstack
Xbias_nstack_0[6] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[6]/vcasc
+ bias_nstack
Xbias_nstack_0[7] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[7]/vcasc
+ bias_nstack
Xbias_nstack_0[8] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[8]/vcasc
+ bias_nstack
Xbias_nstack_0[9] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[9]/vcasc
+ bias_nstack
Xbias_nstack_0[10] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[10]/vcasc
+ bias_nstack
Xbias_nstack_0[11] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[11]/vcasc
+ bias_nstack
Xbias_nstack_0[12] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[12]/vcasc
+ bias_nstack
Xbias_nstack_0[13] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[13]/vcasc
+ bias_nstack
Xbias_nstack_0[14] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[14]/vcasc
+ bias_nstack
Xbias_nstack_0[15] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[15]/vcasc
+ bias_nstack
Xbias_nstack_0[16] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[16]/vcasc
+ bias_nstack
Xbias_nstack_0[17] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[17]/vcasc
+ bias_nstack
Xbias_nstack_0[18] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[18]/vcasc
+ bias_nstack
Xbias_nstack_0[19] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[19]/vcasc
+ bias_nstack
Xbias_nstack_0[20] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[20]/vcasc
+ bias_nstack
Xbias_nstack_0[21] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[21]/vcasc
+ bias_nstack
Xbias_nstack_0[22] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[22]/vcasc
+ bias_nstack
Xbias_nstack_0[23] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[23]/vcasc
+ bias_nstack
Xbias_nstack_0[24] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[24]/vcasc
+ bias_nstack
Xbias_nstack_0[25] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[25]/vcasc
+ bias_nstack
Xbias_nstack_0[26] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[26]/vcasc
+ bias_nstack
Xbias_nstack_0[27] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[27]/vcasc
+ bias_nstack
Xbias_nstack_0[28] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[28]/vcasc
+ bias_nstack
Xbias_nstack_0[29] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[29]/vcasc
+ bias_nstack
Xbias_nstack_0[30] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[30]/vcasc
+ bias_nstack
Xbias_nstack_0[31] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[31]/vcasc
+ bias_nstack
Xbias_nstack_0[32] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[32]/vcasc
+ bias_nstack
Xbias_nstack_0[33] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[33]/vcasc
+ bias_nstack
Xbias_nstack_0[34] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[34]/vcasc
+ bias_nstack
Xbias_nstack_0[35] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[35]/vcasc
+ bias_nstack
Xbias_nstack_0[36] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[36]/vcasc
+ bias_nstack
Xbias_nstack_0[37] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[37]/vcasc
+ bias_nstack
Xbias_nstack_0[38] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[38]/vcasc
+ bias_nstack
Xbias_nstack_0[39] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[39]/vcasc
+ bias_nstack
Xbias_nstack_0[40] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[40]/vcasc
+ bias_nstack
Xbias_nstack_0[41] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[41]/vcasc
+ bias_nstack
Xbias_nstack_0[42] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[43] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[44] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[45] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[46] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[47] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[48] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[49] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[50] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[51] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[52] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[53] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[54] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[55] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[56] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[57] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[58] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[59] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[60] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[61] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[62] bias_pstack_0[62]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[62]/vcasc
+ bias_nstack
Xbias_nstack_0[63] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[63]/vcasc
+ bias_nstack
Xbias_nstack_0[64] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[64]/vcasc
+ bias_nstack
Xbias_nstack_0[65] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[65]/vcasc
+ bias_nstack
Xbias_nstack_0[66] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[66]/vcasc
+ bias_nstack
Xbias_nstack_0[67] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[67]/vcasc
+ bias_nstack
Xbias_nstack_0[68] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[68]/vcasc
+ bias_nstack
Xbias_nstack_0[69] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[69]/vcasc
+ bias_nstack
Xbias_nstack_0[70] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[70]/vcasc
+ bias_nstack
Xbias_nstack_0[71] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[71]/vcasc
+ bias_nstack
Xbias_nstack_0[72] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[72]/vcasc
+ bias_nstack
Xbias_nstack_0[73] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[73]/vcasc
+ bias_nstack
Xbias_nstack_0[74] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[74]/vcasc
+ bias_nstack
Xbias_nstack_0[75] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[75]/vcasc
+ bias_nstack
Xbias_nstack_0[76] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[76]/vcasc
+ bias_nstack
Xbias_nstack_0[77] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[77]/vcasc
+ bias_nstack
Xbias_nstack_0[78] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[78]/vcasc
+ bias_nstack
Xbias_nstack_0[79] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[79]/vcasc
+ bias_nstack
Xbias_nstack_0[80] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[80]/vcasc
+ bias_nstack
Xbias_nstack_0[81] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[81]/vcasc
+ bias_nstack
Xbias_nstack_0[82] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[82]/vcasc
+ bias_nstack
Xbias_nstack_0[83] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[83]/vcasc
+ bias_nstack
Xbias_nstack_0[84] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[84]/vcasc
+ bias_nstack
Xbias_nstack_0[85] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[85]/vcasc
+ bias_nstack
Xbias_nstack_0[86] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[86]/vcasc
+ bias_nstack
Xbias_nstack_0[87] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[87]/vcasc
+ bias_nstack
Xbias_nstack_0[88] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[88]/vcasc
+ bias_nstack
Xbias_nstack_0[89] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[89]/vcasc
+ bias_nstack
Xbias_nstack_0[90] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[90]/vcasc
+ bias_nstack
Xbias_nstack_0[91] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[91]/vcasc
+ bias_nstack
Xbias_nstack_0[92] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[92]/vcasc
+ bias_nstack
Xbias_nstack_0[93] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[93]/vcasc
+ bias_nstack
Xbias_nstack_0[94] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[94]/vcasc
+ bias_nstack
Xbias_nstack_0[95] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[95]/vcasc
+ bias_nstack
Xbias_nstack_0[96] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[96]/vcasc
+ bias_nstack
Xbias_nstack_0[97] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[97]/vcasc
+ bias_nstack
Xbias_nstack_0[98] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[98]/vcasc
+ bias_nstack
Xbias_nstack_0[99] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[99]/vcasc
+ bias_nstack
Xbias_nstack_0[100] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[100]/vcasc
+ bias_nstack
Xbias_nstack_0[101] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[101]/vcasc
+ bias_nstack
Xbias_nstack_0[102] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[102]/vcasc
+ bias_nstack
Xbias_nstack_0[103] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[103]/vcasc
+ bias_nstack
Xbias_nstack_0[104] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[104]/vcasc
+ bias_nstack
Xbias_nstack_0[105] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[105]/vcasc
+ bias_nstack
Xbias_nstack_0[106] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[106]/vcasc
+ bias_nstack
Xbias_nstack_0[107] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[107]/vcasc
+ bias_nstack
Xbias_nstack_0[108] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[108]/vcasc
+ bias_nstack
Xbias_nstack_0[109] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[109]/vcasc
+ bias_nstack
Xbias_nstack_0[110] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[110]/vcasc
+ bias_nstack
Xbias_nstack_0[111] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[111]/vcasc
+ bias_nstack
Xbias_nstack_0[112] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[112]/vcasc
+ bias_nstack
Xbias_nstack_0[113] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[113]/vcasc
+ bias_nstack
Xbias_nstack_0[114] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[114]/vcasc
+ bias_nstack
Xbias_nstack_0[115] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[115]/vcasc
+ bias_nstack
Xbias_nstack_0[116] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[116]/vcasc
+ bias_nstack
Xbias_nstack_0[117] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[117]/vcasc
+ bias_nstack
Xbias_nstack_0[118] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[118]/vcasc
+ bias_nstack
Xbias_nstack_0[119] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[119]/vcasc
+ bias_nstack
Xbias_nstack_0[120] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[120]/vcasc
+ bias_nstack
Xbias_nstack_0[121] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[121]/vcasc
+ bias_nstack
Xbias_nstack_0[122] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[122]/vcasc
+ bias_nstack
Xbias_nstack_0[123] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[123]/vcasc
+ bias_nstack
Xbias_nstack_0[124] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[124]/vcasc
+ bias_nstack
Xbias_nstack_0[125] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[125]/vcasc
+ bias_nstack
Xbias_nstack_0[126] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[126]/vcasc
+ bias_nstack
Xbias_nstack_0[127] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[127]/vcasc
+ bias_nstack
Xbias_nstack_0[128] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[128]/vcasc
+ bias_nstack
Xbias_nstack_0[129] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[129]/vcasc
+ bias_nstack
Xbias_nstack_0[130] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[130]/vcasc
+ bias_nstack
Xbias_nstack_0[131] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[131]/vcasc
+ bias_nstack
Xbias_nstack_0[132] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[132]/vcasc
+ bias_nstack
Xbias_nstack_0[133] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[133]/vcasc
+ bias_nstack
Xbias_nstack_0[134] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[134]/vcasc
+ bias_nstack
Xbias_nstack_0[135] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[135]/vcasc
+ bias_nstack
Xbias_nstack_0[136] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[136]/vcasc
+ bias_nstack
Xbias_nstack_0[137] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[137]/vcasc
+ bias_nstack
Xbias_nstack_0[138] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[138]/vcasc
+ bias_nstack
Xbias_nstack_0[139] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[139]/vcasc
+ bias_nstack
Xbias_nstack_0[140] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[140]/vcasc
+ bias_nstack
Xbias_nstack_0[141] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[141]/vcasc
+ bias_nstack
Xbias_nstack_0[142] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[142]/vcasc
+ bias_nstack
Xbias_nstack_0[143] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[143]/vcasc
+ bias_nstack
Xbias_nstack_0[144] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[144]/vcasc
+ bias_nstack
Xbias_nstack_0[145] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[145]/vcasc
+ bias_nstack
Xbias_nstack_0[146] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[146]/vcasc
+ bias_nstack
Xbias_nstack_0[147] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[147]/vcasc
+ bias_nstack
Xbias_nstack_0[148] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[148]/vcasc
+ bias_nstack
Xbias_nstack_0[149] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[149]/vcasc
+ bias_nstack
Xbias_nstack_0[150] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[150]/vcasc
+ bias_nstack
Xbias_nstack_0[151] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[151]/vcasc
+ bias_nstack
Xbias_nstack_0[152] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[152]/vcasc
+ bias_nstack
Xbias_nstack_0[153] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[153]/vcasc
+ bias_nstack
Xbias_nstack_0[154] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[154]/vcasc
+ bias_nstack
Xbias_nstack_0[155] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[155]/vcasc
+ bias_nstack
Xbias_nstack_0[156] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[156]/vcasc
+ bias_nstack
Xbias_nstack_0[157] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[157]/vcasc
+ bias_nstack
Xbias_nstack_0[158] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[158]/vcasc
+ bias_nstack
Xbias_nstack_0[159] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[159]/vcasc
+ bias_nstack
Xbias_nstack_0[160] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[160]/vcasc
+ bias_nstack
Xbias_nstack_0[161] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[161]/vcasc
+ bias_nstack
Xbias_nstack_0[162] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[162]/vcasc
+ bias_nstack
Xbias_nstack_0[163] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[163]/vcasc
+ bias_nstack
Xbias_nstack_0[164] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[164]/vcasc
+ bias_nstack
Xbias_nstack_0[165] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[165]/vcasc
+ bias_nstack
Xbias_nstack_0[166] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[166]/vcasc
+ bias_nstack
Xbias_nstack_0[167] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[167]/vcasc
+ bias_nstack
Xbias_nstack_0[168] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[168]/vcasc
+ bias_nstack
Xbias_nstack_0[169] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[169]/vcasc
+ bias_nstack
Xbias_nstack_0[170] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[170]/vcasc
+ bias_nstack
Xbias_nstack_0[171] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[171]/vcasc
+ bias_nstack
Xbias_nstack_0[172] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[172]/vcasc
+ bias_nstack
Xbias_nstack_0[173] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[173]/vcasc
+ bias_nstack
Xbias_nstack_0[174] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[174]/vcasc
+ bias_nstack
Xbias_nstack_0[175] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[175]/vcasc
+ bias_nstack
Xbias_nstack_0[176] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[176]/vcasc
+ bias_nstack
Xbias_nstack_0[177] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[177]/vcasc
+ bias_nstack
Xbias_nstack_0[178] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[178]/vcasc
+ bias_nstack
Xbias_nstack_0[179] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[179]/vcasc
+ bias_nstack
Xbias_nstack_0[180] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[180]/vcasc
+ bias_nstack
Xbias_nstack_0[181] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[181]/vcasc
+ bias_nstack
Xbias_nstack_0[182] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[182]/vcasc
+ bias_nstack
Xbias_nstack_0[183] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[183]/vcasc
+ bias_nstack
Xbias_nstack_0[184] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[184]/vcasc
+ bias_nstack
Xbias_nstack_0[185] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[185]/vcasc
+ bias_nstack
Xbias_nstack_0[186] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[186]/vcasc
+ bias_nstack
Xbias_nstack_0[187] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[187]/vcasc
+ bias_nstack
Xbias_nstack_0[188] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[188]/vcasc
+ bias_nstack
Xbias_nstack_0[189] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[189]/vcasc
+ bias_nstack
Xbias_nstack_0[190] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[190]/vcasc
+ bias_nstack
Xbias_nstack_0[191] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[191]/vcasc
+ bias_nstack
Xbias_nstack_0[192] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[192]/vcasc
+ bias_nstack
Xbias_nstack_0[193] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[193]/vcasc
+ bias_nstack
Xbias_nstack_0[194] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[194]/vcasc
+ bias_nstack
Xbias_nstack_0[195] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[195]/vcasc
+ bias_nstack
Xbias_nstack_0[196] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[196]/vcasc
+ bias_nstack
Xbias_nstack_0[197] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[197]/vcasc
+ bias_nstack
Xbias_nstack_0[198] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[198]/vcasc
+ bias_nstack
Xbias_nstack_0[199] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[199]/vcasc
+ bias_nstack
Xbias_nstack_0[200] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[200]/vcasc
+ bias_nstack
Xbias_nstack_0[201] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[201]/vcasc
+ bias_nstack
Xbias_nstack_0[202] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[202]/vcasc
+ bias_nstack
Xbias_nstack_0[203] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[203]/vcasc
+ bias_nstack
Xbias_nstack_0[204] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[204]/vcasc
+ bias_nstack
Xbias_nstack_0[205] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[205]/vcasc
+ bias_nstack
Xbias_nstack_0[206] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[206]/vcasc
+ bias_nstack
Xbias_nstack_0[207] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[207]/vcasc
+ bias_nstack
Xbias_nstack_0[208] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[208]/vcasc
+ bias_nstack
Xbias_nstack_0[209] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[209]/vcasc
+ bias_nstack
Xbias_nstack_0[210] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[210]/vcasc
+ bias_nstack
Xbias_nstack_0[211] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[211]/vcasc
+ bias_nstack
Xbias_nstack_0[212] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[212]/vcasc
+ bias_nstack
Xbias_nstack_0[213] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[213]/vcasc
+ bias_nstack
Xbias_nstack_0[214] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[214]/vcasc
+ bias_nstack
Xbias_nstack_0[215] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[215]/vcasc
+ bias_nstack
Xbias_nstack_0[216] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[216]/vcasc
+ bias_nstack
Xbias_nstack_0[217] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[217]/vcasc
+ bias_nstack
Xbias_nstack_0[218] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[218]/vcasc
+ bias_nstack
Xbias_nstack_0[219] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[219]/vcasc
+ bias_nstack
Xbias_nstack_0[220] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[220]/vcasc
+ bias_nstack
Xbias_nstack_0[221] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[221]/vcasc
+ bias_nstack
Xbias_nstack_0[222] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[222]/vcasc
+ bias_nstack
Xbias_nstack_0[223] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[223]/vcasc
+ bias_nstack
Xbias_nstack_0[224] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[224]/vcasc
+ bias_nstack
Xbias_nstack_0[225] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[225]/vcasc
+ bias_nstack
Xbias_nstack_0[226] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[226]/vcasc
+ bias_nstack
Xbias_nstack_0[227] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[227]/vcasc
+ bias_nstack
Xbias_nstack_0[228] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[228]/vcasc
+ bias_nstack
Xbias_nstack_0[229] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[229]/vcasc
+ bias_nstack
Xbias_nstack_0[230] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[230]/vcasc
+ bias_nstack
Xbias_nstack_0[231] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[231]/vcasc
+ bias_nstack
Xbias_nstack_0[232] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[232]/vcasc
+ bias_nstack
Xbias_nstack_0[233] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[233]/vcasc
+ bias_nstack
Xbias_nstack_0[234] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[234]/vcasc
+ bias_nstack
Xbias_nstack_0[235] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[235]/vcasc
+ bias_nstack
Xbias_nstack_0[236] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[236]/vcasc
+ bias_nstack
Xbias_nstack_0[237] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[237]/vcasc
+ bias_nstack
Xbias_nstack_0[238] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[238]/vcasc
+ bias_nstack
Xbias_nstack_0[239] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[239]/vcasc
+ bias_nstack
Xbias_nstack_0[240] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[240]/vcasc
+ bias_nstack
Xbias_nstack_0[241] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[241]/vcasc
+ bias_nstack
Xbias_nstack_0[242] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[242]/vcasc
+ bias_nstack
Xbias_nstack_0[243] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[243]/vcasc
+ bias_nstack
Xbias_nstack_0[244] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[244]/vcasc
+ bias_nstack
Xbias_nstack_0[245] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[245]/vcasc
+ bias_nstack
Xbias_nstack_0[246] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[246]/vcasc
+ bias_nstack
Xbias_nstack_0[247] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[247]/vcasc
+ bias_nstack
Xbias_nstack_0[248] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[248]/vcasc
+ bias_nstack
Xbias_nstack_0[249] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[249]/vcasc
+ bias_nstack
Xbias_nstack_0[250] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[250]/vcasc
+ bias_nstack
Xbias_nstack_0[251] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[251]/vcasc
+ bias_nstack
Xbias_nstack_0[252] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[252]/vcasc
+ bias_nstack
Xbias_nstack_0[253] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[253]/vcasc
+ bias_nstack
Xbias_nstack_0[254] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[254]/vcasc
+ bias_nstack
Xbias_nstack_0[255] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[255]/vcasc
+ bias_nstack
Xbias_nstack_0[256] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[256]/vcasc
+ bias_nstack
Xbias_nstack_0[257] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[257]/vcasc
+ bias_nstack
Xbias_nstack_0[258] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[258]/vcasc
+ bias_nstack
Xbias_nstack_0[259] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[259]/vcasc
+ bias_nstack
Xbias_nstack_0[260] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[260]/vcasc
+ bias_nstack
Xbias_nstack_0[261] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[261]/vcasc
+ bias_nstack
Xbias_nstack_0[262] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[262]/vcasc
+ bias_nstack
Xbias_nstack_0[263] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[263]/vcasc
+ bias_nstack
Xbias_nstack_0[264] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[264]/vcasc
+ bias_nstack
Xbias_nstack_0[265] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[265]/vcasc
+ bias_nstack
Xbias_nstack_0[266] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[266]/vcasc
+ bias_nstack
Xbias_nstack_0[267] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[267]/vcasc
+ bias_nstack
Xbias_nstack_0[268] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[268]/vcasc
+ bias_nstack
Xbias_nstack_0[269] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[269]/vcasc
+ bias_nstack
Xbias_nstack_0[270] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[270]/vcasc
+ bias_nstack
Xbias_nstack_0[271] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[271]/vcasc
+ bias_nstack
Xbias_nstack_0[272] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[272]/vcasc
+ bias_nstack
Xbias_nstack_0[273] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[273]/vcasc
+ bias_nstack
Xbias_nstack_0[274] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[274]/vcasc
+ bias_nstack
Xbias_nstack_0[275] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[275]/vcasc
+ bias_nstack
Xbias_nstack_0[276] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[276]/vcasc
+ bias_nstack
Xbias_nstack_0[277] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[277]/vcasc
+ bias_nstack
Xbias_nstack_0[278] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[278]/vcasc
+ bias_nstack
Xbias_nstack_0[279] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[279]/vcasc
+ bias_nstack
Xbias_nstack_0[280] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[280]/vcasc
+ bias_nstack
Xbias_nstack_0[281] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[281]/vcasc
+ bias_nstack
Xbias_nstack_0[282] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[282]/vcasc
+ bias_nstack
Xbias_nstack_0[283] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[283]/vcasc
+ bias_nstack
Xbias_nstack_0[284] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[284]/vcasc
+ bias_nstack
Xbias_nstack_0[285] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[285]/vcasc
+ bias_nstack
Xbias_nstack_0[286] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[286]/vcasc
+ bias_nstack
Xbias_nstack_0[287] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[287]/vcasc
+ bias_nstack
Xbias_nstack_0[288] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[288]/vcasc
+ bias_nstack
Xbias_nstack_0[289] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[289]/vcasc
+ bias_nstack
Xbias_nstack_0[290] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[290]/vcasc
+ bias_nstack
Xbias_nstack_0[291] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[291]/vcasc
+ bias_nstack
Xbias_nstack_0[292] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[292]/vcasc
+ bias_nstack
Xbias_nstack_0[293] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[293]/vcasc
+ bias_nstack
Xbias_nstack_0[294] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[294]/vcasc
+ bias_nstack
Xbias_nstack_0[295] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[295]/vcasc
+ bias_nstack
Xbias_nstack_0[296] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[296]/vcasc
+ bias_nstack
Xbias_nstack_0[297] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[297]/vcasc
+ bias_nstack
Xbias_nstack_0[298] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[298]/vcasc
+ bias_nstack
Xbias_nstack_0[299] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[299]/vcasc
+ bias_nstack
Xbias_nstack_0[300] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[300]/vcasc
+ bias_nstack
Xbias_nstack_0[301] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[301]/vcasc
+ bias_nstack
Xbias_nstack_0[302] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[302]/vcasc
+ bias_nstack
Xbias_nstack_0[303] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[303]/vcasc
+ bias_nstack
Xbias_nstack_0[304] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[304]/vcasc
+ bias_nstack
Xbias_nstack_0[305] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[305]/vcasc
+ bias_nstack
Xbias_nstack_0[306] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[306]/vcasc
+ bias_nstack
Xbias_nstack_0[307] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[307]/vcasc
+ bias_nstack
Xbias_nstack_0[308] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[308]/vcasc
+ bias_nstack
Xbias_nstack_0[309] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[309]/vcasc
+ bias_nstack
Xbias_nstack_0[310] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[310]/vcasc
+ bias_nstack
Xbias_nstack_0[311] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[311]/vcasc
+ bias_nstack
Xbias_nstack_0[312] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[312]/vcasc
+ bias_nstack
Xbias_nstack_0[313] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[313]/vcasc
+ bias_nstack
Xbias_nstack_0[314] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[314]/vcasc
+ bias_nstack
Xbias_nstack_0[315] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[315]/vcasc
+ bias_nstack
Xbias_nstack_0[316] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[316]/vcasc
+ bias_nstack
Xbias_nstack_0[317] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[317]/vcasc
+ bias_nstack
Xbias_nstack_0[318] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[318]/vcasc
+ bias_nstack
Xbias_nstack_0[319] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[319]/vcasc
+ bias_nstack
Xbias_nstack_0[320] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[320]/vcasc
+ bias_nstack
Xbias_nstack_0[321] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[321]/vcasc
+ bias_nstack
Xbias_nstack_0[322] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[322]/vcasc
+ bias_nstack
Xbias_nstack_0[323] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[323]/vcasc
+ bias_nstack
Xbias_nstack_0[324] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[324]/vcasc
+ bias_nstack
Xbias_nstack_0[325] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[325]/vcasc
+ bias_nstack
Xbias_nstack_0[326] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[326]/vcasc
+ bias_nstack
Xbias_nstack_0[327] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[327]/vcasc
+ bias_nstack
Xbias_nstack_0[328] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[328]/vcasc
+ bias_nstack
Xbias_nstack_0[329] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[329]/vcasc
+ bias_nstack
Xbias_nstack_0[330] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[330]/vcasc
+ bias_nstack
Xbias_nstack_0[331] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[331]/vcasc
+ bias_nstack
Xbias_nstack_0[332] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[332]/vcasc
+ bias_nstack
Xbias_nstack_0[333] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[333]/vcasc
+ bias_nstack
Xbias_nstack_0[334] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[334]/vcasc
+ bias_nstack
Xbias_nstack_0[335] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[335]/vcasc
+ bias_nstack
Xbias_nstack_0[336] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[336]/vcasc
+ bias_nstack
Xbias_nstack_0[337] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[337]/vcasc
+ bias_nstack
Xbias_nstack_0[338] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[338]/vcasc
+ bias_nstack
Xbias_nstack_0[339] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[339]/vcasc
+ bias_nstack
Xbias_nstack_0[340] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[340]/vcasc
+ bias_nstack
Xbias_nstack_0[341] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[341]/vcasc
+ bias_nstack
Xbias_nstack_0[342] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[342]/vcasc
+ bias_nstack
Xbias_nstack_0[343] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[343]/vcasc
+ bias_nstack
Xbias_nstack_0[344] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[344]/vcasc
+ bias_nstack
Xbias_nstack_0[345] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[345]/vcasc
+ bias_nstack
Xbias_nstack_0[346] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[346]/vcasc
+ bias_nstack
Xbias_nstack_0[347] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[347]/vcasc
+ bias_nstack
Xbias_nstack_0[348] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[348]/vcasc
+ bias_nstack
Xbias_nstack_0[349] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[349]/vcasc
+ bias_nstack
Xbias_nstack_0[350] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[350]/vcasc
+ bias_nstack
Xbias_nstack_0[351] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[351]/vcasc
+ bias_nstack
Xbias_nstack_0[352] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[352]/vcasc
+ bias_nstack
Xbias_nstack_0[353] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[353]/vcasc
+ bias_nstack
Xbias_nstack_0[354] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[354]/vcasc
+ bias_nstack
Xbias_nstack_0[355] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[355]/vcasc
+ bias_nstack
Xbias_nstack_0[356] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[356]/vcasc
+ bias_nstack
Xbias_nstack_0[357] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[357]/vcasc
+ bias_nstack
Xbias_nstack_0[358] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[358]/vcasc
+ bias_nstack
Xbias_nstack_0[359] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[359]/vcasc
+ bias_nstack
Xbias_nstack_0[360] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[360]/vcasc
+ bias_nstack
Xbias_nstack_0[361] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[361]/vcasc
+ bias_nstack
Xbias_nstack_0[362] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[362]/vcasc
+ bias_nstack
Xbias_nstack_0[363] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[363]/vcasc
+ bias_nstack
Xbias_nstack_0[364] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[364]/vcasc
+ bias_nstack
Xbias_nstack_0[365] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[365]/vcasc
+ bias_nstack
Xbias_nstack_0[366] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[366]/vcasc
+ bias_nstack
Xbias_nstack_0[367] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[367]/vcasc
+ bias_nstack
Xbias_nstack_0[368] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[368]/vcasc
+ bias_nstack
Xbias_nstack_0[369] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[369]/vcasc
+ bias_nstack
Xbias_nstack_0[370] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[370]/vcasc
+ bias_nstack
Xbias_nstack_0[371] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[371]/vcasc
+ bias_nstack
Xbias_nstack_0[372] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[372]/vcasc
+ bias_nstack
Xbias_nstack_0[373] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[373]/vcasc
+ bias_nstack
Xbias_nstack_0[374] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[374]/vcasc
+ bias_nstack
Xbias_nstack_0[375] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[375]/vcasc
+ bias_nstack
Xbias_nstack_0[376] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[376]/vcasc
+ bias_nstack
Xbias_nstack_0[377] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[377]/vcasc
+ bias_nstack
Xbias_nstack_0[378] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[378]/vcasc
+ bias_nstack
Xbias_nstack_0[379] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[379]/vcasc
+ bias_nstack
Xbias_nstack_0[380] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[380]/vcasc
+ bias_nstack
Xbias_nstack_0[381] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[381]/vcasc
+ bias_nstack
Xbias_nstack_0[382] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[382]/vcasc
+ bias_nstack
Xbias_nstack_0[383] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[383]/vcasc
+ bias_nstack
Xbias_nstack_0[384] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[384]/vcasc
+ bias_nstack
Xbias_nstack_0[385] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[385]/vcasc
+ bias_nstack
Xbias_nstack_0[386] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[386]/vcasc
+ bias_nstack
Xbias_nstack_0[387] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[387]/vcasc
+ bias_nstack
Xbias_nstack_0[388] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[388]/vcasc
+ bias_nstack
Xbias_nstack_0[389] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[389]/vcasc
+ bias_nstack
Xbias_nstack_0[390] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[390]/vcasc
+ bias_nstack
Xbias_nstack_0[391] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[391]/vcasc
+ bias_nstack
Xbias_nstack_0[392] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[392]/vcasc
+ bias_nstack
Xbias_nstack_0[393] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[393]/vcasc
+ bias_nstack
Xbias_nstack_0[394] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[394]/vcasc
+ bias_nstack
Xbias_nstack_0[395] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[395]/vcasc
+ bias_nstack
Xbias_nstack_0[396] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[396]/vcasc
+ bias_nstack
Xbias_nstack_0[397] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[397]/vcasc
+ bias_nstack
Xbias_nstack_0[398] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[398]/vcasc
+ bias_nstack
Xbias_nstack_0[399] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[399]/vcasc
+ bias_nstack
Xbias_nstack_0[400] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[400]/vcasc
+ bias_nstack
Xbias_nstack_0[401] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[401]/vcasc
+ bias_nstack
Xbias_nstack_0[402] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[402]/vcasc
+ bias_nstack
Xbias_nstack_0[403] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[403]/vcasc
+ bias_nstack
Xbias_nstack_0[404] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[404]/vcasc
+ bias_nstack
Xbias_nstack_0[405] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[405]/vcasc
+ bias_nstack
Xbias_nstack_0[406] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[406]/vcasc
+ bias_nstack
Xbias_nstack_0[407] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[407]/vcasc
+ bias_nstack
Xbias_nstack_0[408] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[408]/vcasc
+ bias_nstack
Xbias_nstack_0[409] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[409]/vcasc
+ bias_nstack
Xbias_nstack_0[410] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[410]/vcasc
+ bias_nstack
Xbias_nstack_0[411] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[411]/vcasc
+ bias_nstack
Xbias_nstack_0[412] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[412]/vcasc
+ bias_nstack
Xbias_nstack_0[413] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[413]/vcasc
+ bias_nstack
Xbias_nstack_0[414] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[414]/vcasc
+ bias_nstack
Xbias_nstack_0[415] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[415]/vcasc
+ bias_nstack
Xbias_nstack_0[416] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[416]/vcasc
+ bias_nstack
Xbias_nstack_0[417] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[417]/vcasc
+ bias_nstack
Xbias_nstack_0[418] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[418]/vcasc
+ bias_nstack
Xbias_nstack_0[419] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[419]/vcasc
+ bias_nstack
Xbias_nstack_0[420] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[420]/vcasc
+ bias_nstack
Xbias_nstack_0[421] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[421]/vcasc
+ bias_nstack
Xbias_nstack_0[422] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[422]/vcasc
+ bias_nstack
Xbias_nstack_0[423] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[423]/vcasc
+ bias_nstack
Xbias_nstack_0[424] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[424]/vcasc
+ bias_nstack
Xbias_nstack_0[425] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[425]/vcasc
+ bias_nstack
Xbias_nstack_0[426] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[426]/vcasc
+ bias_nstack
Xbias_nstack_0[427] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[427]/vcasc
+ bias_nstack
Xbias_nstack_0[428] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[428]/vcasc
+ bias_nstack
Xbias_nstack_0[429] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[429]/vcasc
+ bias_nstack
Xbias_nstack_0[430] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[430]/vcasc
+ bias_nstack
Xbias_nstack_0[431] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[431]/vcasc
+ bias_nstack
Xbias_nstack_0[432] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[432]/vcasc
+ bias_nstack
Xbias_nstack_0[433] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[433]/vcasc
+ bias_nstack
Xbias_nstack_0[434] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[434]/vcasc
+ bias_nstack
Xbias_nstack_0[435] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[435]/vcasc
+ bias_nstack
Xbias_nstack_0[436] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[436]/vcasc
+ bias_nstack
Xbias_nstack_0[437] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[437]/vcasc
+ bias_nstack
Xbias_nstack_0[438] snk_test1 ena_test1 bias_nstack_0[9]/nbias avss bias_nstack_0[438]/vcasc
+ bias_nstack
Xbias_nstack_0[439] snk_test1 ena_test1 bias_nstack_0[9]/nbias avss bias_nstack_0[439]/vcasc
+ bias_nstack
XXR2 m1_6353_1231# m1_11831_n5169# m1_2369_1231# m1_10005_1231# m1_9175_n5169# m1_4527_n5169#
+ m1_5855_n5169# m1_5357_1231# m1_10835_n5169# m1_10337_1231# m1_8179_n5169# m1_5025_1231#
+ m1_2037_1231# m1_5523_n5169# m1_12163_n5169# ref_in m1_8345_1231# m1_211_n5169#
+ m1_11333_1231# m1_6353_1231# m1_2369_1231# m1_7183_n5169# m1_11167_n5169# m1_12495_n5169#
+ m1_1207_n5169# m1_8013_1231# m1_11001_1231# m1_10171_n5169# m1_11499_n5169# m1_11333_1231#
+ m1_n121_n5169# m1_6851_n5169# m1_2701_1231# m1_4029_1231# m1_n287_1231# m1_8345_1231#
+ m1_5855_n5169# m1_2203_n5169# m1_10669_1231# m1_875_n5169# m1_6021_1231# m1_10503_n5169#
+ m1_3199_n5169# m1_4361_1231# m1_1373_1231# m1_45_1231# bias_pstack_0[9]/pcasc m1_12163_n5169#
+ m1_1871_n5169# m1_9009_1231# m1_9507_n5169# m1_6685_1231# m1_4195_n5169# m1_11001_1231#
+ m1_11167_n5169# m1_5025_1231# m1_8511_n5169# m1_12329_1231# m1_4693_1231# m1_2867_n5169#
+ m1_1705_1231# m1_1539_n5169# m1_9341_1231# m1_5191_n5169# m1_11665_1231# m1_6519_n5169#
+ m1_6685_1231# m1_10171_n5169# m1_3863_n5169# m1_2535_n5169# m1_2037_1231# m1_7515_n5169#
+ m1_8677_1231# m1_9175_n5169# m1_6851_n5169# m1_3531_n5169# m1_1705_1231# m1_9009_1231#
+ m1_11997_1231# m1_11831_n5169# m1_4859_n5169# m1_n453_n5169# m1_3697_1231# m1_1871_n5169#
+ m1_8677_1231# m1_709_1231# m1_8179_n5169# m1_11665_1231# m1_7349_1231# m1_4527_n5169#
+ m1_543_n5169# m1_10835_n5169# m1_5523_n5169# m1_4029_1231# m1_2867_n5169# m1_1041_1231#
+ m1_7183_n5169# m1_5689_1231# m1_9673_1231# m1_12495_n5169# m1_6187_n5169# m1_211_n5169#
+ avss m1_9839_n5169# m1_3697_1231# m1_709_1231# m1_7017_1231# m1_10005_1231# m1_3863_n5169#
+ m1_n121_n5169# m1_4361_1231# m1_1373_1231# m1_11499_n5169# m1_5689_1231# m1_9673_1231#
+ m1_1207_n5169# bias_nstack_0[61]/itail m1_4859_n5169# m1_8843_n5169# m1_875_n5169#
+ m1_n453_n5169# m1_7017_1231# m1_10503_n5169# m1_1041_1231# m1_2203_n5169# m1_3033_1231#
+ m1_7847_n5169# m1_9507_n5169# m1_2701_1231# m1_9341_1231# m1_6187_n5169# m1_n287_1231#
+ m1_8013_1231# m1_12329_1231# m1_543_n5169# m1_3199_n5169# m1_6021_1231# m1_3365_1231#
+ m1_1539_n5169# m1_377_1231# bias_pstack_0[9]/pcasc m1_8511_n5169# m1_10669_1231#
+ m1_11997_1231# m1_9839_n5169# m1_4195_n5169# m1_2535_n5169# m1_45_1231# m1_5191_n5169#
+ m1_7515_n5169# m1_5357_1231# m1_8843_n5169# m1_6519_n5169# m1_3033_1231# m1_4693_1231#
+ m1_377_1231# m1_7349_1231# m1_7847_n5169# m1_10337_1231# m1_3531_n5169# m1_3365_1231#
+ sky130_fd_pr__res_high_po_0p35_P35QVK
Xbias_pstack_0[0] bias_pstack_0[9]/pcasc enb_test0 src_test0 bias_pstack_0[0]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[1] bias_pstack_0[9]/pcasc enb_test0 src_test0 bias_pstack_0[1]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[2] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[2]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[3] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[3]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[4] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[4]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[5] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[5]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[6] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[6]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[7] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[7]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[8] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[8]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[9] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[9]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[10] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[10]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[11] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[11]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[12] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[12]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[13] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[13]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[14] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[14]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[15] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[15]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[16] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[16]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[17] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[17]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[18] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[18]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[19] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[19]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[20] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[20]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[21] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[21]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[22] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[22]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[23] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[23]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[24] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[24]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[25] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[25]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[26] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[26]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[27] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[27]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[28] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[28]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[29] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[29]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[30] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[30]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[31] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[31]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[32] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[32]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[33] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[33]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[34] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[34]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[35] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[35]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[36] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[36]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[37] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[37]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[38] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[38]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[39] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[39]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[40] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[40]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[41] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[41]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[42] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[42]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[43] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[43]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[44] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[44]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[45] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[45]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[46] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[46]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[47] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[47]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[48] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[48]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[49] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[49]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[50] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[50]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[51] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[51]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[52] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[52]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[53] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[53]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[54] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[54]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[55] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[55]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[56] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[56]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[57] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[57]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[58] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[58]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[59] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[59]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[60] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[60]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[61] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[61]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[62] bias_pstack_0[9]/pcasc enb bias_pstack_0[62]/itail bias_pstack_0[9]/pbias
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[63] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[63]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[64] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[64]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[65] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[65]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[66] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[66]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[67] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[67]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[68] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[68]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[69] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[69]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[70] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[70]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[71] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[71]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[72] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[72]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[73] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[73]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[74] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[74]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[75] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[75]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[76] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[76]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[77] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[77]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[78] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[78]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[79] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[79]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[80] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[80]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[81] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[81]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[82] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[82]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[83] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[83]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[84] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[84]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[85] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[85]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[86] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[86]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[87] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[87]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[88] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[88]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[89] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[89]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[90] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[90]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[91] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[91]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[92] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[92]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[93] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[93]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[94] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[94]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[95] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[95]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[96] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[96]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[97] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[97]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[98] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[98]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[99] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[99]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[100] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[100]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[101] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[101]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[102] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[102]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[103] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[103]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[104] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[104]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[105] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[105]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[106] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[106]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[107] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[107]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[108] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[108]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[109] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[109]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[110] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[110]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[111] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[111]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[112] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[112]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[113] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[113]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[114] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[114]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[115] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[115]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[116] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[116]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[117] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[117]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[118] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[118]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[119] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[119]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[120] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[120]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[121] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[121]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[122] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[122]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[123] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[123]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[124] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[124]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[125] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[125]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[126] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[126]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[127] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[127]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[128] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[128]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[129] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[129]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[130] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[130]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[131] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[131]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[132] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[132]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[133] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[133]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[134] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[134]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[135] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[135]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[136] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[136]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[137] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[137]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[138] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[138]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[139] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[139]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[140] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[140]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[141] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[141]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[142] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[142]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[143] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[143]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[144] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[144]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[145] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[145]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[146] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[146]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[147] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[147]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[148] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[148]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[149] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[149]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[150] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[150]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[151] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[151]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[152] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[152]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[153] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[153]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[154] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[154]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[155] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[155]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[156] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[156]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[157] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[157]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[158] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[158]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[159] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[159]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[160] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[160]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[161] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[161]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[162] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[162]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[163] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[163]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[164] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[164]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[165] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[165]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[166] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[166]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[167] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[167]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[168] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[168]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[169] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[169]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[170] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[170]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[171] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[171]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[172] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[172]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[173] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[173]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[174] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[174]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[175] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[175]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[176] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[176]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[177] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[177]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[178] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[178]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[179] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[179]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[180] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[180]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[181] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[181]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[182] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[182]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[183] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[183]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[184] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[184]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[185] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[185]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[186] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[186]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[187] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[187]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[188] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[188]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[189] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[189]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[190] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[190]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[191] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[191]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[192] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[192]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[193] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[193]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[194] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[194]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[195] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[195]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[196] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[196]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[197] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[197]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[198] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[198]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[199] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[199]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[200] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[200]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[201] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[201]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[202] bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[202]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[203] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[203]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[204] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[204]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[205] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[205]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[206] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[206]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[207] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[207]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[208] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[208]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[209] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[209]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[210] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[210]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[211] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[211]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[212] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[212]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[213] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[213]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[214] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[214]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[215] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[215]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[216] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[216]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[217] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[217]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[218] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[218]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[219] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[219]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[220] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[220]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[221] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[221]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[222] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[222]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[223] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[223]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[224] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[224]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[225] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[225]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[226] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[226]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[227] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[227]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[228] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[228]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[229] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[229]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[230] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[230]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[231] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[231]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[232] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[232]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[233] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[233]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[234] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[234]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[235] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[235]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[236] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[236]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[237] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[237]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[238] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[238]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[239] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[239]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[240] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[240]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[241] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[241]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[242] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[242]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[243] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[243]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[244] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[244]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[245] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[245]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[246] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[246]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[247] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[247]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[248] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[248]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[249] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[249]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[250] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[250]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[251] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[251]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[252] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[252]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[253] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[253]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[254] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[254]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[255] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[255]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[256] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[256]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[257] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[257]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[258] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[258]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[259] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[259]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[260] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[260]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[261] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[261]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[262] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[262]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[263] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[263]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[264] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[264]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[265] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[265]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[266] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[266]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[267] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[267]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[268] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[268]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[269] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[269]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[270] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[270]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[271] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[271]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[272] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[272]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[273] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[273]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[274] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[274]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[275] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[275]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[276] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[276]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[277] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[277]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[278] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[278]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[279] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[279]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[280] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[280]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[281] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[281]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[282] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[282]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[283] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[283]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[284] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[284]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[285] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[285]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[286] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[286]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[287] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[287]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[288] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[288]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[289] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[289]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[290] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[290]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[291] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[291]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[292] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[292]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[293] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[293]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[294] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[294]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[295] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[295]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[296] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[296]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[297] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[297]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[298] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[298]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[299] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[299]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[300] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[300]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[301] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[301]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[302] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[302]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[303] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[303]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[304] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[304]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[305] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[305]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[306] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[306]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[307] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[307]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[308] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[308]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[309] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[309]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[310] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[310]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[311] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[311]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[312] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[312]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[313] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[313]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[314] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[314]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[315] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[315]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[316] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[316]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[317] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[317]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[318] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[318]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[319] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[319]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[320] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[320]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[321] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[321]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[322] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[322]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[323] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[323]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[324] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[324]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[325] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[325]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[326] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[326]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[327] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[327]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[328] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[328]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[329] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[329]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[330] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[330]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[331] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[331]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[332] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[332]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[333] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[333]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[334] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[334]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[335] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[335]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[336] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[336]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[337] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[337]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[338] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[338]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[339] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[339]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[340] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[340]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[341] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[341]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[342] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[342]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[343] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[343]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[344] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[344]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[345] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[345]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[346] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[346]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[347] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[347]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[348] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[348]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[349] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[349]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[350] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[350]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[351] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[351]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[352] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[352]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[353] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[353]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[354] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[354]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[355] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[355]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[356] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[356]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[357] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[357]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[358] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[358]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[359] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[359]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[360] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[360]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[361] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[361]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[362] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[362]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[363] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[363]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[364] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[364]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[365] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[365]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[366] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[366]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[367] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[367]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[368] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[368]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[369] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[369]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[370] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[370]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[371] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[371]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[372] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[372]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[373] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[373]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[374] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[374]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[375] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[375]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[376] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[376]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[377] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[377]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[378] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[378]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[379] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[379]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[380] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[380]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[381] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[381]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[382] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[382]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[383] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[383]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[384] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[384]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[385] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[385]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[386] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[386]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[387] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[387]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[388] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[388]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[389] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[389]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[390] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[390]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[391] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[391]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[392] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[392]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[393] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[393]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[394] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[394]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[395] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[395]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[396] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[396]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[397] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[397]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[398] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[398]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[399] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[399]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[400] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[400]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[401] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[401]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[402] bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[402]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[403] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[403]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[404] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[404]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[405] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[405]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[406] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[406]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[407] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[407]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[408] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[408]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[409] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[409]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[410] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[410]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[411] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[411]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[412] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[412]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[413] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[413]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[414] bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[414]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[415] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[415]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[416] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[416]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[417] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[417]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[418] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[418]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[419] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[419]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[420] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[420]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[421] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[421]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[422] bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[422]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[423] bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[423]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[424] bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[424]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[425] bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[425]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[426] bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[426]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[427] bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[427]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[428] bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[428]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[429] bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[429]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[430] bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[430]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[431] bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[431]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[432] bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[432]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[433] bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[433]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[434] bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[434]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[435] bias_pstack_0[9]/pcasc enb_100 src_100 bias_pstack_0[435]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[436] bias_pstack_0[9]/pcasc enb_100 src_100 bias_pstack_0[436]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[437] bias_pstack_0[9]/pcasc enb_50 src_50 bias_pstack_0[437]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[438] bias_pstack_0[9]/pcasc enb_test1 src_test1 bias_pstack_0[438]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[439] bias_pstack_0[9]/pcasc enb_test1 src_test1 bias_pstack_0[439]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WQT6C6 a_1235_n700# a_3447_n700# a_5659_n700#
+ a_n287_n788# a_761_n700# a_n4079_n788# a_819_n788# a_2657_n700# a_4869_n700# a_5185_n700#
+ a_n1077_n788# a_n3289_n788# a_1867_n700# a_2183_n700# a_345_n788# a_4395_n700# a_n29_n700#
+ a_n2499_n788# a_1393_n700# a_n919_n788# a_6607_n700# a_977_n788# a_n5027_n788# a_3605_n700#
+ a_5817_n700# a_n445_n788# a_3189_n788# a_n187_n700# a_6133_n700# a_n1709_n788# a_n2025_n788#
+ a_n4237_n788# a_2815_n700# a_n6449_n788# a_3131_n700# a_5343_n700# a_2399_n788#
+ a_n1235_n788# a_n3447_n788# a_n5659_n788# a_n3189_n700# a_2341_n700# a_4553_n700#
+ a_503_n788# a_6765_n700# a_n2657_n788# a_n4869_n788# a_n5185_n788# a_n2399_n700#
+ a_1551_n700# a_3763_n700# a_5975_n700# a_1609_n788# a_6291_n700# a_n1867_n788# a_6349_n788#
+ a_n819_n700# a_4137_n788# a_n2183_n788# a_n4395_n788# a_2973_n700# a_n603_n788#
+ a_3347_n788# a_1135_n788# a_n7124_n700# a_n345_n700# a_5559_n788# a_n1393_n788#
+ a_n1609_n700# a_n6607_n788# a_661_n788# a_n6349_n700# a_n4137_n700# a_5501_n700#
+ a_4769_n788# a_2557_n788# a_5085_n788# a_n3605_n788# a_n5817_n788# a_n3347_n700#
+ a_n1135_n700# a_n6133_n788# a_n5559_n700# a_4711_n700# a_6923_n700# a_3979_n788#
+ a_1767_n788# a_n977_n700# a_4295_n788# a_2083_n788# a_n2815_n788# a_n3131_n788#
+ a_n5343_n788# a_n4769_n700# a_n2557_n700# a_3921_n700# a_n5085_n700# a_1293_n788#
+ a_n761_n788# a_6507_n788# a_n2341_n788# a_n3979_n700# a_n1767_n700# a_n4553_n788#
+ a_n6765_n788# a_n4295_n700# a_n2083_n700# a_5717_n788# a_3505_n788# a_6033_n788#
+ a_n503_n700# a_n1551_n788# a_n3763_n788# a_n5975_n788# a_n1293_n700# a_129_n700#
+ a_n6291_n788# a_n6507_n700# a_2715_n788# a_4927_n788# a_3031_n788# a_n2973_n788#
+ a_5243_n788# a_n5717_n700# a_n3505_n700# a_n6033_n700# a_1925_n788# a_4453_n788#
+ a_2241_n788# a_6665_n788# a_n2715_n700# a_n5501_n788# a_n4927_n700# a_n3031_n700#
+ a_n5243_n700# a_1451_n788# a_5875_n788# a_n661_n700# a_3663_n788# a_6191_n788# a_287_n700#
+ a_n4711_n788# a_n1925_n700# a_n6923_n788# a_n4453_n700# a_n2241_n700# a_n6665_n700#
+ a_2873_n788# a_n3921_n788# a_n1451_n700# a_n5875_n700# a_n3663_n700# a_n6191_n700#
+ a_5401_n788# a_n2873_n700# a_6823_n788# a_4611_n788# a_919_n700# a_n5401_n700# a_3821_n788#
+ a_445_n700# a_n6823_n700# a_n4611_n700# a_n3821_n700# a_4079_n700# a_1077_n700#
+ a_3289_n700# a_29_n788# a_2499_n700# a_n6981_n700# a_n129_n788# a_603_n700# a_187_n788#
+ a_5027_n700# a_1709_n700# a_2025_n700# a_4237_n700# a_6449_n700#
X0 a_n6349_n700# a_n6449_n788# a_n6507_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X1 a_n5875_n700# a_n5975_n788# a_n6033_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X2 a_n3505_n700# a_n3605_n788# a_n3663_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X3 a_3605_n700# a_3505_n788# a_3447_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X4 a_5975_n700# a_5875_n788# a_5817_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X5 a_6449_n700# a_6349_n788# a_6291_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X6 a_n6191_n700# a_n6291_n788# a_n6349_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X7 a_n977_n700# a_n1077_n788# a_n1135_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X8 a_6291_n700# a_6191_n788# a_6133_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X9 a_n503_n700# a_n603_n788# a_n661_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X10 a_1077_n700# a_977_n788# a_919_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X11 a_n5401_n700# a_n5501_n788# a_n5559_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X12 a_n2557_n700# a_n2657_n788# a_n2715_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X13 a_2657_n700# a_2557_n788# a_2499_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X14 a_5501_n700# a_5401_n788# a_5343_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X15 a_n4927_n700# a_n5027_n788# a_n5085_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X16 a_n4453_n700# a_n4553_n788# a_n4611_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X17 a_n29_n700# a_n129_n788# a_n187_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X18 a_603_n700# a_503_n788# a_445_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X19 a_4553_n700# a_4453_n788# a_4395_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X20 a_n6507_n700# a_n6607_n788# a_n6665_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X21 a_6607_n700# a_6507_n788# a_6449_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X22 a_n3979_n700# a_n4079_n788# a_n4137_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X23 a_n1135_n700# a_n1235_n788# a_n1293_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X24 a_1235_n700# a_1135_n788# a_1077_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X25 a_5659_n700# a_5559_n788# a_5501_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X26 a_n5559_n700# a_n5659_n788# a_n5717_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X27 a_n2715_n700# a_n2815_n788# a_n2873_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X28 a_2815_n700# a_2715_n788# a_2657_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X29 a_n3031_n700# a_n3131_n788# a_n3189_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X30 a_3131_n700# a_3031_n788# a_2973_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X31 a_n4611_n700# a_n4711_n788# a_n4769_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X32 a_n1767_n700# a_n1867_n788# a_n1925_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X33 a_1867_n700# a_1767_n788# a_1709_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X34 a_4711_n700# a_4611_n788# a_4553_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X35 a_2183_n700# a_2083_n788# a_2025_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X36 a_n2083_n700# a_n2183_n788# a_n2241_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X37 a_n4137_n700# a_n4237_n788# a_n4295_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X38 a_n3663_n700# a_n3763_n788# a_n3821_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X39 a_3763_n700# a_3663_n788# a_3605_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X40 a_4237_n700# a_4137_n788# a_4079_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X41 a_n819_n700# a_n919_n788# a_n977_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X42 a_n5717_n700# a_n5817_n788# a_n5875_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X43 a_n661_n700# a_n761_n788# a_n819_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X44 a_5817_n700# a_5717_n788# a_5659_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X45 a_n6033_n700# a_n6133_n788# a_n6191_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X46 a_n3189_n700# a_n3289_n788# a_n3347_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X47 a_3289_n700# a_3189_n788# a_3131_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X48 a_6133_n700# a_6033_n788# a_5975_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X49 a_n4769_n700# a_n4869_n788# a_n4927_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X50 a_919_n700# a_819_n788# a_761_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X51 a_2025_n700# a_1925_n788# a_1867_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X52 a_4869_n700# a_4769_n788# a_4711_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X53 a_n5085_n700# a_n5185_n788# a_n5243_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X54 a_n187_n700# a_n287_n788# a_n345_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X55 a_761_n700# a_661_n788# a_603_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X56 a_5185_n700# a_5085_n788# a_5027_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X57 a_n2241_n700# a_n2341_n788# a_n2399_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X58 a_2341_n700# a_2241_n788# a_2183_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X59 a_n6665_n700# a_n6765_n788# a_n6823_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X60 a_n3821_n700# a_n3921_n788# a_n3979_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X61 a_287_n700# a_187_n788# a_129_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X62 a_3921_n700# a_3821_n788# a_3763_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X63 a_6765_n700# a_6665_n788# a_6607_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X64 a_n1293_n700# a_n1393_n788# a_n1451_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X65 a_1393_n700# a_1293_n788# a_1235_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X66 a_n3347_n700# a_n3447_n788# a_n3505_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X67 a_n2873_n700# a_n2973_n788# a_n3031_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X68 a_2973_n700# a_2873_n788# a_2815_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X69 a_3447_n700# a_3347_n788# a_3289_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X70 a_5027_n700# a_4927_n788# a_4869_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X71 a_n345_n700# a_n445_n788# a_n503_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X72 a_2499_n700# a_2399_n788# a_2341_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X73 a_5343_n700# a_5243_n788# a_5185_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X74 a_n5243_n700# a_n5343_n788# a_n5401_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X75 a_n2399_n700# a_n2499_n788# a_n2557_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X76 a_n6823_n700# a_n6923_n788# a_n6981_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X77 a_n1609_n700# a_n1709_n788# a_n1767_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X78 a_129_n700# a_29_n788# a_n29_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X79 a_1709_n700# a_1609_n788# a_1551_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X80 a_4079_n700# a_3979_n788# a_3921_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X81 a_6923_n700# a_6823_n788# a_6765_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X82 a_n4295_n700# a_n4395_n788# a_n4453_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X83 a_n1925_n700# a_n2025_n788# a_n2083_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X84 a_n1451_n700# a_n1551_n788# a_n1609_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X85 a_445_n700# a_345_n788# a_287_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X86 a_1551_n700# a_1451_n788# a_1393_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X87 a_4395_n700# a_4295_n788# a_4237_n700# a_n7124_n700# sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7WGKBW a_5875_n1597# a_5343_n1500# a_n761_n1597#
+ a_3131_n1500# a_5817_n1500# a_3663_n1597# a_187_n1597# a_129_n1500# a_3605_n1500#
+ a_1451_n1597# a_1925_n1597# a_n2399_n1500# a_n6133_n1597# a_5185_n1500# a_661_n1597#
+ a_n6607_n1597# a_5659_n1500# a_603_n1500# a_3447_n1500# a_3979_n1597# a_1293_n1597#
+ a_n2873_n1500# a_1767_n1597# a_1235_n1500# a_1709_n1500# a_n6449_n1597# a_3921_n1500#
+ a_977_n1597# a_445_n1500# a_n4237_n1597# a_919_n1500# a_3289_n1500# a_n2025_n1597#
+ a_6033_n1597# a_1077_n1500# a_6507_n1597# a_n6923_n1597# a_5975_n1500# a_n5401_n1500#
+ a_n4711_n1597# a_287_n1500# a_3763_n1500# a_n4079_n1597# a_1551_n1500# a_n6291_n1597#
+ a_6349_n1597# a_n6765_n1597# a_761_n1500# a_n5243_n1500# a_n29_n1500# a_4137_n1597#
+ a_n4553_n1597# a_n5717_n1500# a_n3031_n1500# a_n2341_n1597# a_1393_n1500# a_n3505_n1500#
+ a_n2815_n1597# a_6823_n1597# a_1867_n1500# a_4611_n1597# a_n5085_n1500# a_n4395_n1597#
+ a_n5559_n1500# a_6191_n1597# a_n2183_n1597# a_n4869_n1597# a_n3347_n1500# a_6665_n1597#
+ a_6133_n1500# a_n2657_n1597# a_n1135_n1500# a_6607_n1500# a_4453_n1597# a_n1609_n1500#
+ a_4927_n1597# a_n503_n1500# a_2241_n1597# a_n3821_n1500# a_2715_n1597# a_n3189_n1500#
+ a_n2499_n1597# a_6449_n1500# a_4295_n1597# a_n5875_n1500# a_4237_n1500# a_4769_n1597#
+ a_2083_n1597# a_n345_n1500# a_n3663_n1500# a_2025_n1500# a_2557_n1597# a_n2973_n1597#
+ a_n819_n1500# a_n1451_n1500# a_6923_n1500# a_n1925_n1500# a_4711_n1500# a_29_n1597#
+ a_n5027_n1597# a_4079_n1500# a_n187_n1500# a_2399_n1597# a_6291_n1500# a_n3979_n1500#
+ a_n1293_n1500# a_6765_n1500# a_n1767_n1500# a_n5501_n1597# a_4553_n1500# a_n661_n1500#
+ a_2341_n1500# a_2873_n1597# a_2815_n1500# a_n6033_n1500# a_n5343_n1597# a_n6507_n1500#
+ a_4395_n1500# a_n3131_n1597# a_n5817_n1597# a_n977_n1500# a_2183_n1500# a_4869_n1500#
+ a_n3605_n1597# a_2657_n1500# a_5401_n1597# a_n5185_n1597# a_n6349_n1500# a_n5659_n1597#
+ a_n129_n1597# a_n4137_n1500# a_n3447_n1597# a_2499_n1500# a_5243_n1597# a_n1235_n1597#
+ a_n1709_n1597# a_n6823_n1500# a_5717_n1597# a_3031_n1597# a_n603_n1597# a_n4611_n1500#
+ a_3505_n1597# a_n3921_n1597# a_2973_n1500# a_n3289_n1597# a_n1077_n1597# a_n6191_n1500#
+ a_5085_n1597# w_n7017_n1600# a_n6665_n1500# a_5027_n1500# a_5559_n1597# a_503_n1597#
+ a_n5975_n1597# a_n445_n1597# a_n4453_n1500# a_3347_n1597# a_n3763_n1597# a_n919_n1597#
+ a_n4927_n1500# a_n2241_n1500# a_1135_n1597# a_n1551_n1597# a_n2715_n1500# a_1609_n1597#
+ a_5501_n1500# a_3821_n1597# a_345_n1597# a_n287_n1597# a_n4295_n1500# a_3189_n1597#
+ a_819_n1597# a_n4769_n1500# a_n2083_n1500# a_n1393_n1597# a_n6981_n1500# a_n2557_n1500#
+ a_n1867_n1597#
X0 a_n6033_n1500# a_n6133_n1597# a_n6191_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X1 a_n819_n1500# a_n919_n1597# a_n977_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X2 a_n6191_n1500# a_n6291_n1597# a_n6349_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X3 a_n977_n1500# a_n1077_n1597# a_n1135_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X4 a_2973_n1500# a_2873_n1597# a_2815_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X5 a_n6507_n1500# a_n6607_n1597# a_n6665_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X6 a_1235_n1500# a_1135_n1597# a_1077_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X7 a_1393_n1500# a_1293_n1597# a_1235_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X8 a_4079_n1500# a_3979_n1597# a_3921_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X9 a_n6665_n1500# a_n6765_n1597# a_n6823_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X10 a_603_n1500# a_503_n1597# a_445_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X11 a_1709_n1500# a_1609_n1597# a_1551_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X12 a_n4927_n1500# a_n5027_n1597# a_n5085_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X13 a_761_n1500# a_661_n1597# a_603_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X14 a_6923_n1500# a_6823_n1597# a_6765_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=0.5
X15 a_n5085_n1500# a_n5185_n1597# a_n5243_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X16 a_n4453_n1500# a_n4553_n1597# a_n4611_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X17 a_n3821_n1500# a_n3921_n1597# a_n3979_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X18 a_1867_n1500# a_1767_n1597# a_1709_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X19 a_2499_n1500# a_2399_n1597# a_2341_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X20 a_4711_n1500# a_4611_n1597# a_4553_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X21 a_5343_n1500# a_5243_n1597# a_5185_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X22 a_n2241_n1500# a_n2341_n1597# a_n2399_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X23 a_n5559_n1500# a_n5659_n1597# a_n5717_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X24 a_3131_n1500# a_3031_n1597# a_2973_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X25 a_n503_n1500# a_n603_n1597# a_n661_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X26 a_5817_n1500# a_5717_n1597# a_5659_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X27 a_6449_n1500# a_6349_n1597# a_6291_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X28 a_n3347_n1500# a_n3447_n1597# a_n3505_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X29 a_n2715_n1500# a_n2815_n1597# a_n2873_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X30 a_287_n1500# a_187_n1597# a_129_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X31 a_5975_n1500# a_5875_n1597# a_5817_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X32 a_n3979_n1500# a_n4079_n1597# a_n4137_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X33 a_n2873_n1500# a_n2973_n1597# a_n3031_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X34 a_n661_n1500# a_n761_n1597# a_n819_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X35 a_3605_n1500# a_3505_n1597# a_3447_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X36 a_4237_n1500# a_4137_n1597# a_4079_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X37 a_n1135_n1500# a_n1235_n1597# a_n1293_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X38 a_3763_n1500# a_3663_n1597# a_3605_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X39 a_4395_n1500# a_4295_n1597# a_4237_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X40 a_n1293_n1500# a_n1393_n1597# a_n1451_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X41 a_n6823_n1500# a_n6923_n1597# a_n6981_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=0.5
X42 a_n1609_n1500# a_n1709_n1597# a_n1767_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X43 a_n29_n1500# a_n129_n1597# a_n187_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X44 a_1551_n1500# a_1451_n1597# a_1393_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X45 a_2183_n1500# a_2083_n1597# a_2025_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X46 a_4869_n1500# a_4769_n1597# a_4711_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X47 a_n1767_n1500# a_n1867_n1597# a_n1925_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X48 a_n187_n1500# a_n287_n1597# a_n345_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X49 a_n4611_n1500# a_n4711_n1597# a_n4769_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X50 a_n2399_n1500# a_n2499_n1597# a_n2557_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X51 a_2025_n1500# a_1925_n1597# a_1867_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X52 a_n5243_n1500# a_n5343_n1597# a_n5401_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X53 a_2657_n1500# a_2557_n1597# a_2499_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X54 a_3289_n1500# a_3189_n1597# a_3131_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X55 a_5501_n1500# a_5401_n1597# a_5343_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X56 a_6133_n1500# a_6033_n1597# a_5975_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X57 a_n5717_n1500# a_n5817_n1597# a_n5875_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X58 a_n3031_n1500# a_n3131_n1597# a_n3189_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X59 a_129_n1500# a_29_n1597# a_n29_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X60 a_n6349_n1500# a_n6449_n1597# a_n6507_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X61 a_6291_n1500# a_6191_n1597# a_6133_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X62 a_n5875_n1500# a_n5975_n1597# a_n6033_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X63 a_445_n1500# a_345_n1597# a_287_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X64 a_6607_n1500# a_6507_n1597# a_6449_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X65 a_n4137_n1500# a_n4237_n1597# a_n4295_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X66 a_n3505_n1500# a_n3605_n1597# a_n3663_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X67 a_6765_n1500# a_6665_n1597# a_6607_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X68 a_n3663_n1500# a_n3763_n1597# a_n3821_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X69 a_n4295_n1500# a_n4395_n1597# a_n4453_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X70 a_n1925_n1500# a_n2025_n1597# a_n2083_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X71 a_919_n1500# a_819_n1597# a_761_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X72 a_3921_n1500# a_3821_n1597# a_3763_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X73 a_4553_n1500# a_4453_n1597# a_4395_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X74 a_n1451_n1500# a_n1551_n1597# a_n1609_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X75 a_1077_n1500# a_977_n1597# a_919_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X76 a_5185_n1500# a_5085_n1597# a_5027_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X77 a_n4769_n1500# a_n4869_n1597# a_n4927_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X78 a_n2083_n1500# a_n2183_n1597# a_n2241_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X79 a_2341_n1500# a_2241_n1597# a_2183_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X80 a_5027_n1500# a_4927_n1597# a_4869_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X81 a_5659_n1500# a_5559_n1597# a_5501_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X82 a_n2557_n1500# a_n2657_n1597# a_n2715_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X83 a_n345_n1500# a_n445_n1597# a_n503_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X84 a_n5401_n1500# a_n5501_n1597# a_n5559_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X85 a_n3189_n1500# a_n3289_n1597# a_n3347_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X86 a_2815_n1500# a_2715_n1597# a_2657_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
X87 a_3447_n1500# a_3347_n1597# a_3289_n1500# w_n7017_n1600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3BH9ZH a_n345_n200# a_129_n200# a_287_n200# a_428_n196#
+ a_29_n288# a_n129_n288# a_187_n288# a_n287_n288# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n288# a_n29_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n288# a_n187_n200# a_428_n196# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RTDP6L a_n29_n400# w_n381_n500# a_n187_n400#
+ a_n345_n400# a_29_n497# a_n129_n497# a_187_n497# a_129_n400# a_n287_n497# a_287_n400#
X0 a_n29_n400# a_n129_n497# a_n187_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n187_n400# a_n287_n497# a_n345_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2 a_287_n400# a_187_n497# a_129_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X3 a_129_n400# a_29_n497# a_n29_n400# w_n381_n500# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt gate_drive in_m in_p out vdd vss vsub
Xxm1 vss vss vss li_n2466_n1927# out li_n5626_n1927# li_n2466_n1927# out out out li_n2466_n1927#
+ li_n5626_n1927# vss vss li_n2466_n1927# vss vss li_n2466_n1927# out li_n2466_n1927#
+ vss li_n2466_n1927# li_n5626_n1927# out out li_n2466_n1927# li_n2466_n1927# out
+ out li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# vss li_n6574_n1927# vss vss
+ li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# li_n5626_n1927# vss out out li_n2466_n1927#
+ out li_n5626_n1927# li_n5626_n1927# li_n5626_n1927# out vss vss vss li_n2466_n1927#
+ vss li_n2466_n1927# li_n2466_n1927# out li_n2466_n1927# li_n2466_n1927# li_n5626_n1927#
+ out li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# vss vss li_n2466_n1927# li_n2466_n1927#
+ vss li_n6574_n1927# li_n2466_n1927# vss vss out li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# li_n5626_n1927# li_n6574_n1927# li_n2466_n1927# out li_n6574_n1927#
+ li_n2466_n1927# vss vss li_n2466_n1927# li_n2466_n1927# vss li_n2466_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n5626_n1927# li_n5626_n1927# vss vss out vss li_n2466_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# out li_n5626_n1927#
+ li_n7839_364# li_n2466_n1927# out li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ out li_n2466_n1927# li_n5626_n1927# li_n6574_n1927# vss out li_n6574_n1927# li_n5626_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# li_n2466_n1927#
+ vss vss vss li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# vss li_n2466_n1927# li_n2466_n1927# vss li_n5626_n1927# vss li_n7839_364#
+ vss vss vss li_n2466_n1927# li_n5626_n1927# out li_n5626_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# vss li_n2466_n1927# li_n2466_n1927# vss vss li_n2466_n1927#
+ out li_n6574_n1927# li_n2466_n1927# vss vss out out li_n2466_n1927# vss vss li_n2466_n1927#
+ vss li_n2466_n1927# vss out out out out sky130_fd_pr__nfet_g5v0d10v5_WQT6C6
Xxm2 li_n2466_n1927# vdd li_n2466_n1927# vdd out li_n2466_n1927# li_n2466_n1927# out
+ out li_n2466_n1927# li_n2466_n1927# out li_n6574_n1927# out li_n2466_n1927# li_n6574_n1927#
+ vdd vdd vdd li_n2466_n1927# li_n2466_n1927# vdd li_n2466_n1927# vdd out li_n6574_n1927#
+ out li_n2466_n1927# out li_n5626_n1927# vdd out li_n2466_n1927# li_n2466_n1927#
+ out li_n2466_n1927# li_n7839_364# vdd vdd li_n5626_n1927# vdd vdd li_n5626_n1927#
+ vdd li_n6574_n1927# li_n2466_n1927# li_n7839_364# out li_n2466_n1927# vdd li_n2466_n1927#
+ li_n5626_n1927# vdd li_n2466_n1927# li_n2466_n1927# out vdd li_n5626_n1927# li_n2466_n1927#
+ vdd li_n2466_n1927# vdd li_n5626_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# li_n2466_n1927# out li_n5626_n1927# out vdd li_n2466_n1927#
+ vdd li_n2466_n1927# out li_n2466_n1927# vdd li_n2466_n1927# vdd li_n2466_n1927#
+ out li_n2466_n1927# li_n5626_n1927# out li_n2466_n1927# li_n2466_n1927# vdd li_n2466_n1927#
+ out li_n2466_n1927# li_n5626_n1927# out out vdd vdd vdd li_n2466_n1927# li_n5626_n1927#
+ vdd out li_n2466_n1927# vdd li_n2466_n1927# vdd out out li_n5626_n1927# out vdd
+ out li_n2466_n1927# vdd vdd li_n5626_n1927# li_n5626_n1927# vdd li_n5626_n1927#
+ li_n6574_n1927# vdd vdd out li_n5626_n1927# out li_n2466_n1927# li_n5626_n1927#
+ vdd li_n5626_n1927# li_n2466_n1927# vdd li_n5626_n1927# vdd li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# li_n6574_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n5626_n1927# out li_n5626_n1927# li_n2466_n1927#
+ li_n5626_n1927# li_n2466_n1927# vdd vdd vdd li_n2466_n1927# li_n2466_n1927# li_n6574_n1927#
+ li_n2466_n1927# vdd li_n2466_n1927# li_n5626_n1927# li_n2466_n1927# li_n2466_n1927#
+ vdd li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# out li_n2466_n1927#
+ li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927# li_n2466_n1927#
+ vdd out li_n2466_n1927# vdd vdd li_n2466_n1927# sky130_fd_pr__pfet_g5v0d10v5_7WGKBW
Xxm3 vss li_n7839_364# vss vss in_m in_p in_m in_p vss li_n7529_279# sky130_fd_pr__nfet_g5v0d10v5_3BH9ZH
Xxm4 vdd vdd li_n7529_279# vdd li_n7529_279# li_n7839_364# li_n7529_279# li_n7839_364#
+ li_n7839_364# vdd sky130_fd_pr__pfet_g5v0d10v5_RTDP6L
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt pmos_waffle_48x48 dw_n11050_n11060# w_n10844_n10854# a_n50_n50# a_112_3350#
+ a_112_1150#
X0 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X5 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X6 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X7 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X8 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X9 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X10 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X11 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X12 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X13 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X14 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X15 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X16 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X17 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X18 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X19 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X20 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X21 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X22 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X23 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X24 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X25 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X26 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X27 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X28 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X29 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X30 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X31 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X32 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X33 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X34 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X35 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X36 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X37 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X38 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X39 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X40 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X41 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X42 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X43 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X44 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X45 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X46 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X47 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X48 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X49 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X50 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X51 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X52 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X53 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X54 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X55 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X56 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X57 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X58 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X59 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X60 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X61 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X62 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X63 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X64 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X65 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X66 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X67 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X68 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X69 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X70 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X71 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X72 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X73 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X74 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X75 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X76 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X77 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X78 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X79 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X80 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X81 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X82 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X83 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X84 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X85 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X86 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X87 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X88 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X89 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X90 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X91 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X92 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X93 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X94 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X95 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X96 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X97 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X98 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X99 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X100 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X101 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X103 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X104 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X105 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X106 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X109 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X111 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X113 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X114 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X115 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X116 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X118 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X119 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X120 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X122 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X123 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X125 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X126 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X128 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X129 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X130 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X131 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X132 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X133 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X136 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X137 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X138 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X139 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X140 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X141 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X142 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X143 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X144 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X147 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X148 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X149 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X150 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X151 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X152 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X153 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X154 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X155 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X156 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X157 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X158 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X159 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X160 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X165 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X166 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X167 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X168 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X169 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X171 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X173 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X175 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X176 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X177 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X178 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X179 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X180 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X181 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X182 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X185 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X186 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X187 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X188 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X189 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X190 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X191 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X192 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X193 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X194 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X195 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X196 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X199 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X200 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X201 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X202 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X205 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X207 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X208 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X209 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X210 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X211 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X212 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X213 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X214 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X215 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X216 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X217 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X218 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X219 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X221 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X222 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X224 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X226 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X227 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X228 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X229 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X230 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X231 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X232 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X233 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X235 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X236 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X237 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X238 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X239 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X241 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X243 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X246 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X247 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X248 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X250 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X251 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X252 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X253 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X254 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X255 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X257 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X259 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X260 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X261 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X262 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X263 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X265 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X266 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X267 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X268 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X269 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X270 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X271 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X276 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X278 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X279 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X285 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X286 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X288 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X289 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X290 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X291 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X292 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X293 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X294 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X295 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X296 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X297 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X298 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X299 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X300 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X303 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X305 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X306 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X308 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X310 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X311 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X313 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X314 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X315 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X316 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X320 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X321 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X324 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X325 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X327 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X328 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X329 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X330 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X332 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X334 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X335 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X336 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X337 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X339 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X340 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X341 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X342 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X343 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X344 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X345 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X346 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X347 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X349 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X351 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X352 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X353 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X354 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X356 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X357 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X359 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X360 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X361 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X362 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X363 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X364 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X365 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X366 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X367 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X368 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X369 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X370 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X371 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X373 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X374 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X375 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X376 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X377 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X378 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X381 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X383 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X384 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X386 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X387 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X388 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X389 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X390 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X393 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X394 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X395 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X398 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X399 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X402 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X403 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X404 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X405 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X406 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X407 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X408 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X410 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X411 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X413 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X414 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X415 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X419 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X421 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X422 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X423 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X424 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X425 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X426 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X427 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X431 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X432 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X434 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X435 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X436 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X438 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X440 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X441 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X442 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X443 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X444 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X445 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X446 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X447 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X448 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X451 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X453 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X455 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X457 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X458 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X459 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X460 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X461 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X462 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X463 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X466 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X467 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X468 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X470 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X471 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X474 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X476 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X479 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X480 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X481 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X482 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X483 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X484 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X485 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X486 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X487 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X488 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X489 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X490 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X492 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X493 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X494 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X496 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X499 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X501 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X502 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X503 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X504 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X507 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X509 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X510 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X511 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X512 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X513 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X514 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X515 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X516 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X517 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X518 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X519 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X521 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X522 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X523 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X524 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X525 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X526 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X527 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X528 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X529 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X530 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X531 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X532 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X533 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X534 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X535 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X536 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X537 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X538 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X539 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X540 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X541 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X542 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X543 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X544 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X545 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X546 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X547 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X548 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X549 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X551 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X552 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X553 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X554 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X555 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X556 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X557 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X558 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X559 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X560 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X561 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X562 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X563 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X564 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X565 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X566 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X567 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X569 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X570 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X571 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X572 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X573 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X574 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X575 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X576 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X577 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X578 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X579 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X581 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X582 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X583 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X584 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X585 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X586 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X587 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X588 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X589 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X591 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X592 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X594 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X595 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X596 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X597 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X598 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X599 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X600 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X601 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X602 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X603 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X604 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X605 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X606 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X607 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X608 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X609 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X610 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X611 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X612 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X613 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X614 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X616 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X617 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X619 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X620 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X621 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X622 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X623 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X624 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X625 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X626 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X627 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X628 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X630 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X631 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X632 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X633 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X634 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X635 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X636 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X637 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X638 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X639 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X640 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X641 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X642 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X644 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X645 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X646 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33125 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X647 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X649 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X650 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X652 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X653 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X654 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X655 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X656 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X657 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X658 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X659 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X660 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X661 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X663 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X664 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X665 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X666 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X668 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X669 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X670 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X672 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X673 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X674 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X675 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X676 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X678 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X679 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X680 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X681 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X682 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X683 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X684 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X685 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X686 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X688 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X689 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X690 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X692 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X693 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X694 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X695 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X696 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X697 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X699 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X700 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X701 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X702 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X704 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X705 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X706 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X707 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X708 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X709 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X710 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X711 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X712 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X713 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X714 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X715 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X717 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X718 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X719 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X720 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X721 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X722 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X725 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X727 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X728 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X729 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X731 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X733 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X736 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X737 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X738 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X739 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X740 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X741 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X742 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X743 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X745 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X746 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X747 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X748 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X749 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X751 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X752 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X753 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X754 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X755 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X756 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X757 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X758 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X759 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X760 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X761 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X762 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X763 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X764 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X765 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X768 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X769 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X770 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X771 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X772 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X773 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X774 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X775 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X776 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X777 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X778 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X779 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X781 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X783 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X784 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X785 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X786 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X787 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X788 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X789 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X790 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X791 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X792 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X793 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X794 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X795 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X797 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X799 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X800 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X801 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X802 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X803 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X804 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X805 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X806 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X807 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X809 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X810 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X812 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X814 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X815 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X816 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X817 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X818 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X819 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X820 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X821 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X822 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X823 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X824 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X825 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X826 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X827 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X828 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X829 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X830 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X831 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X833 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X834 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X835 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X836 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X837 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X838 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X839 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X841 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X842 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X843 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X844 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X845 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X846 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X847 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X848 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X849 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X850 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X851 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X852 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X853 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X854 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X855 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X856 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X857 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X858 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X859 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X860 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X861 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X862 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X863 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X864 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X865 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X866 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X867 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X868 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X869 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X870 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X871 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X872 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X873 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X876 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X878 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X879 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X881 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X882 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X883 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X884 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X885 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X886 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X887 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X888 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X889 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X890 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X891 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X892 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X893 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X894 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X895 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X897 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X898 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X899 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X900 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X901 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X903 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X904 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X905 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X906 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X908 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X909 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X910 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X912 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X914 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X915 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X916 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X917 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X918 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X919 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X921 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X922 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X923 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X926 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X927 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X928 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X930 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X931 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X932 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X934 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X935 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X936 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X938 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X939 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X940 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X941 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X942 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X943 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X944 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X945 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X946 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X947 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X948 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X949 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X950 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X951 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X952 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X953 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X954 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X955 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X956 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X957 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X958 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X959 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X960 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X961 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X962 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X964 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X965 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X966 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X967 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X968 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X970 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X971 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X972 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X973 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X974 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X975 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X977 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X978 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X979 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X980 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X981 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X982 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X983 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X984 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X985 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X986 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X987 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X988 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X989 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X990 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X994 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X995 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X996 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X997 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X998 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X999 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1000 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1001 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1003 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1004 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1005 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1007 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1008 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1009 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1010 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1011 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1012 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1013 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1014 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1015 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1016 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1017 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1018 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1020 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1021 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1022 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1023 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1024 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1026 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1027 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1028 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1030 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1031 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1032 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1034 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1035 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1036 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1037 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1038 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1039 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1040 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1041 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1042 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1044 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1045 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1046 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1047 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1048 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1049 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1050 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1051 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1052 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1053 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1054 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1055 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1056 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1057 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1058 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1059 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1060 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1061 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1062 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1063 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1064 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1065 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1066 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1067 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1068 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1069 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1070 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1071 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1072 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1073 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1074 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1075 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1076 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1077 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1078 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1079 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1081 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1082 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1083 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1084 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1085 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1086 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1087 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1088 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1089 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1090 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1091 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1093 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1095 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1096 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1097 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1098 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1100 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1101 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1103 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1104 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1105 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1106 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1109 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1111 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1113 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1114 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1115 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1116 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1118 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1119 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1120 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1122 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1123 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1125 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1126 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1128 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1129 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1130 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1131 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1132 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1133 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1137 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1138 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1139 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1140 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1141 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1142 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1143 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1144 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1145 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1146 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1147 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1148 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1149 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1150 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1153 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1154 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1155 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1156 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1157 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1158 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1159 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1161 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1162 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1165 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1166 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1167 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1168 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1169 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1173 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1175 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1176 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1177 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1178 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1179 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1180 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1181 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1182 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1185 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1186 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1187 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1189 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1190 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1191 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1192 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1193 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1194 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1195 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1196 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1199 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1200 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1201 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1202 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1205 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1207 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1208 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1209 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1210 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1211 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1212 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1214 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1215 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1216 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1217 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1218 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1219 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1221 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1222 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1224 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1225 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1226 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1227 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1228 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1229 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1230 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1231 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1232 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1233 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1235 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1236 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1237 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1238 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1239 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1241 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1243 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1245 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1246 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1247 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1248 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1250 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1251 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1252 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1254 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1255 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1257 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1259 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1260 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1262 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1263 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1265 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1266 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1267 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1269 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1270 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1271 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1272 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1276 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1277 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1278 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1279 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1282 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1286 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1288 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1289 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1290 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1291 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1292 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1293 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1294 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1295 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1296 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1298 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1299 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1300 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1303 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1306 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1308 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1310 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1311 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1314 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1315 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1316 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1320 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1321 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1324 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1325 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1327 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1328 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1329 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1330 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1331 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1332 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1334 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1335 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1336 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1337 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1339 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1340 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1341 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1342 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1343 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1344 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1345 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1347 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1349 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1351 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1352 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1353 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1354 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1356 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1358 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1360 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1361 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1362 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1363 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1364 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1365 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1367 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1368 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1369 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1370 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1371 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1372 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1373 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1374 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1375 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1376 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1377 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1378 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1381 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1383 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1384 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1386 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1387 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1389 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1392 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1393 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1394 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1395 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1402 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1403 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1404 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1405 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1406 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1408 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1409 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1410 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1411 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1413 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1414 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1415 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1416 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1418 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1419 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1421 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1422 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1424 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1425 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1426 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1427 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1431 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1432 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1434 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1436 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1438 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1440 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1441 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1442 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1443 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1444 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1445 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1446 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1447 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1448 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1451 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1453 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1455 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1457 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1458 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1459 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1460 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1461 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1462 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1463 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1464 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1465 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1466 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1467 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1468 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1469 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1470 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1471 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1474 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1475 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1476 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1479 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1480 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1481 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1482 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1483 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1484 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1485 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1486 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1487 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1488 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1489 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1490 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1492 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1493 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1494 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1496 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1497 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1499 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1500 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1503 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1504 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1507 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1509 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1510 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1511 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1512 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1513 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1514 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1515 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1516 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1517 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1518 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1519 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1521 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1522 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1523 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1524 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1525 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1526 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1527 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1528 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1529 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1530 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1531 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1532 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1533 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1534 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1535 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1536 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1537 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1538 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1539 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1540 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1541 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1542 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1543 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1544 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1545 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1546 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1547 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1548 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1549 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1551 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1552 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1553 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1554 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1555 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1556 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1557 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1558 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1559 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1560 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1561 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1562 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1563 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1564 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1565 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1566 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1567 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1569 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1570 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1571 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1572 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1573 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1574 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1575 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1576 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1577 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1578 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1579 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1581 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1582 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1583 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1584 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1585 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1586 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1587 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1588 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1589 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1591 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1592 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1594 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1595 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1596 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1597 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1598 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1599 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1600 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1601 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1602 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1603 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1604 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1605 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1606 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1607 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1608 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1609 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1610 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1611 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1612 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1613 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1614 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1616 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1617 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1619 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1620 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1621 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1622 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1623 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1624 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1625 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1626 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1627 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1628 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1630 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1631 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1632 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1633 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1634 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1635 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1636 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1637 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1638 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1639 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1640 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1641 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1642 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1644 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1645 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1646 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1647 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1649 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1650 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1652 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1653 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1654 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1655 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1656 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1657 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1658 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1659 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1660 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1661 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1663 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1664 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1665 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1666 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1668 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1669 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1670 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1672 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1673 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1674 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1675 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1676 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1678 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1679 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1680 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1681 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1682 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1683 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1684 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1685 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1686 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1688 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1689 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1690 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1692 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1693 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1694 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1695 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1696 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1697 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1699 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1700 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1701 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1702 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1704 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1705 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1706 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1707 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1708 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1709 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1710 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1711 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1712 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1713 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1714 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1715 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1717 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1718 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1719 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1720 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1721 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1722 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1725 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1727 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1728 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1729 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1731 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1733 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1736 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1737 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1738 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1739 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1740 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1741 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1742 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1743 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1745 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1746 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1747 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1748 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1749 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1751 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1752 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1753 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1754 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1755 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1756 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1757 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1758 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1759 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1760 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1761 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1762 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1763 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1764 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1765 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1768 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1769 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1770 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1771 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1772 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1773 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1774 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1775 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1776 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1777 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1778 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1779 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1781 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1783 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1784 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1785 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1786 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1787 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1788 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1789 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1790 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1791 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1792 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1793 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1794 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1795 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1797 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1799 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1800 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1801 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1802 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1803 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1804 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1805 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1806 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1807 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1809 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1810 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1812 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1814 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1815 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1816 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1817 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1818 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1819 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1820 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1821 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1822 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1823 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1824 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1825 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1826 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1827 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1828 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1829 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1830 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1831 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1833 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1834 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1835 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1836 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1837 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1838 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1839 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1841 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1842 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1843 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1844 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1845 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1846 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1847 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1848 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1849 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1850 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1851 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1852 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1853 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1854 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1855 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1856 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1857 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1858 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1859 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1860 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1861 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1862 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1863 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1864 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1865 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1866 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1867 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1868 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1869 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1870 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1871 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1872 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1873 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1876 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1878 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1879 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1881 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1882 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1883 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1884 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1885 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1886 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1887 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1888 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1889 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1890 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1891 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1892 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1893 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1894 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1895 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1897 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1898 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1899 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1900 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1901 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X1902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1903 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1904 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1905 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1906 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1908 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1909 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1910 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1912 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1914 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1915 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1916 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1917 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1918 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1919 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1921 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1922 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X1923 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1926 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1927 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1928 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1930 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1931 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1932 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1934 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1935 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1936 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1938 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1939 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1940 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1941 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1942 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1943 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1944 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1945 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1946 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1947 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1948 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1949 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1950 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1951 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1952 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1953 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1954 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1955 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1956 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1957 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1958 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1959 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1960 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1961 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1962 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1964 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1965 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1966 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1967 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1968 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1970 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1971 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1972 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1973 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1974 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1975 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X1976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1977 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1978 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1979 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X1980 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.33125 ps=9.38 w=4.38 l=0.5
X1981 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1982 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1983 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1984 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1985 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1986 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1987 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1988 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1989 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1990 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X1991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1994 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X1995 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1996 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1997 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X1998 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X1999 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2000 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2001 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2003 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2004 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2005 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2007 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2008 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2009 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2010 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2011 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2012 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2013 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2014 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2015 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2016 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2017 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2018 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2020 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2021 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2022 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2023 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2024 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2026 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2027 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2028 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2030 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2031 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2032 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2034 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2035 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2036 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2037 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2038 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2039 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2040 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2041 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2042 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2044 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2045 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2046 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2047 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2048 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2049 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2050 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2051 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2052 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2053 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2054 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2055 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2056 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2057 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2058 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2059 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2060 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2061 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2062 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2063 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2064 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2065 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2066 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2067 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2068 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2069 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2070 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2071 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2072 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2073 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2074 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2075 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2076 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2077 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2078 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2079 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2081 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2082 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2083 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2084 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2085 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2086 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2087 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2088 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2089 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2090 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2091 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2093 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2095 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2096 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2097 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2098 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2100 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2101 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2103 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2104 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2105 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2106 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2109 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2111 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2113 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2114 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2115 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2116 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2118 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2119 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2120 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2122 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2123 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2124 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2125 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2126 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2128 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2129 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2130 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2131 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2132 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2133 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2137 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2138 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2139 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2140 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2141 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2142 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2143 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2144 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2147 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2148 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2149 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2150 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2153 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2154 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2155 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2156 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2157 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2158 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2159 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2165 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2166 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2167 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2168 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2169 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2173 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2175 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2176 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2177 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2178 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2179 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2180 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2181 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2182 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2184 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2185 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2186 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2187 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2189 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2190 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2191 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2192 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2193 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2194 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2195 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2196 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2197 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2199 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2200 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2201 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2202 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2205 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2207 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2208 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2209 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2210 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2211 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2212 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2214 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2215 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2216 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2217 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2218 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2219 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2220 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2221 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2222 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2224 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2226 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2227 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2228 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2229 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2230 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2231 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2232 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2233 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2235 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2236 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2237 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2238 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2239 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2241 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2243 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2246 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2247 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2248 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2250 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2251 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2252 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2254 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2255 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2257 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2258 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2259 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2260 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2262 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2263 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2264 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2265 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2266 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2267 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2269 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2270 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2271 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2276 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2278 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2279 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2281 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2286 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2287 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2288 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2289 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2290 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2291 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2292 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2293 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2294 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2295 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2296 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2298 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2299 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2300 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2303 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2306 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2308 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2310 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2311 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2314 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2315 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2316 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2318 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2320 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2321 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2322 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2324 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2325 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2327 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2328 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2329 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2330 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2332 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2334 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2335 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2336 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2337 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2339 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2340 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2341 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2342 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2343 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2344 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2345 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2347 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2349 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2351 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2352 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2353 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2354 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2356 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2360 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2361 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2362 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2363 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2364 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2365 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2367 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2368 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2369 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2370 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2371 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2373 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2374 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2375 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2376 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2377 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2378 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2381 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2383 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2384 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2386 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2387 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2389 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2391 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33125 pd=9.38 as=6.2285 ps=16.31 w=4.38 l=0.5
X2393 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2394 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2395 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2402 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2403 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2404 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2405 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2406 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2408 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2410 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2411 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2413 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2414 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2415 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2419 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2421 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2422 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2424 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2425 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2426 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2427 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2430 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2431 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2432 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2434 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2436 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2438 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2440 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2441 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2442 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2443 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2444 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2445 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2446 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2447 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2448 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2450 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2451 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2453 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2455 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2457 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2458 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2459 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2460 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2461 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2462 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2463 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2466 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2467 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2468 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2470 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2471 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2472 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2473 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2474 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2476 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2479 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2480 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2481 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2482 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2483 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2484 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2485 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2486 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2487 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2488 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2489 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2490 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2492 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2493 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2494 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2496 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2499 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2503 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2504 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2507 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2509 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2510 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2511 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2512 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2513 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2514 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2515 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2516 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2517 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2518 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2519 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2521 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2522 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2523 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2524 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2525 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2526 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2527 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2528 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2529 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2530 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2531 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2532 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2533 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2534 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2535 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2536 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2537 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2538 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2539 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2540 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2541 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2542 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2543 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2544 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2545 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2546 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2547 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2548 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2549 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2551 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2552 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2553 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2554 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2555 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2556 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2557 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2558 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2559 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2560 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2561 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2562 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2563 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2564 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2565 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2566 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2567 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2569 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2570 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2571 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2572 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2573 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2574 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2575 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2576 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2577 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2578 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2579 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2581 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2582 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2583 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2584 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2585 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2586 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2587 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2588 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2589 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2591 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2592 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2594 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2595 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2596 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2597 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2598 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2599 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2600 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2601 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2602 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2603 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2604 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2605 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2606 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2607 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2608 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2609 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X2610 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2611 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2612 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2613 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2614 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2616 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2617 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2619 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2620 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2621 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2622 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X2623 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2624 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2625 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2626 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2627 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2628 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2630 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2631 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2632 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2633 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2634 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2635 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2636 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2637 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2638 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2639 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2640 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2641 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2642 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2644 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2645 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2646 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2647 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2649 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2650 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2652 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2653 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2654 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2655 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2656 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2657 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2658 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2659 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2660 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2661 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2663 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2664 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2665 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2666 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2668 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2669 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2670 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2672 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2673 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2674 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2675 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2676 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2678 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2679 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2680 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2681 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2682 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2683 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2684 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2685 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2686 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2688 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2689 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2690 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2692 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2693 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2694 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2695 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2696 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2697 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2699 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2700 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2701 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2702 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2704 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2705 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2706 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2707 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2708 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2709 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2710 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2711 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2712 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2713 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2714 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2715 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2717 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2718 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2719 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2720 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2721 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2722 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2725 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2727 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2728 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2729 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2731 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2733 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2736 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2737 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2738 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2739 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2740 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2741 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2742 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2743 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2745 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2746 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2747 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2748 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2749 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2751 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2752 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2753 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2754 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2755 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2756 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2757 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2758 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2759 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2760 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2761 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2762 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2763 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2764 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2765 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2768 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2769 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2770 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2771 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2772 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2773 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2774 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2775 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2776 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2777 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2778 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2779 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2781 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2783 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2784 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2785 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2786 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2787 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2788 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2789 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2790 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2791 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2792 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2793 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2794 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2795 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2797 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2799 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2800 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2801 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2802 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2803 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2804 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2805 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2806 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2807 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2809 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2810 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2812 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2814 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2815 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2816 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2817 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2818 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2819 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2820 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2821 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2822 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2823 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2824 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2825 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2826 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2827 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2828 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2829 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2830 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2831 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2833 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2834 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2835 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2836 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2837 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2838 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2839 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2841 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2842 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2843 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2844 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2845 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2846 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2847 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2848 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2849 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2850 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2851 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2852 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2853 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2854 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2855 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2856 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2857 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2858 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2859 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2860 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2861 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2862 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2863 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2864 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2865 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2866 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2867 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2868 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2869 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2870 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2871 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2872 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2873 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2876 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2878 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2879 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2881 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2882 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2883 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2884 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2885 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2886 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2887 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2888 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2889 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2890 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2891 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2892 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2893 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2894 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2895 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2897 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2898 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2899 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2900 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2901 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2903 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2904 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2905 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2906 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2908 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2909 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2910 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2912 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2914 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2915 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2916 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2917 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2918 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2919 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2921 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2922 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2923 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2926 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2927 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2928 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X2929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2930 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2931 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2932 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2934 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2935 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2936 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2938 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2939 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2940 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2941 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2942 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2943 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=1.33125 ps=9.38 w=4.38 l=0.5
X2944 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2945 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2946 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2947 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2948 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2949 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2950 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2951 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2952 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2953 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2954 dw_n11050_n11060# a_n50_n50# a_112_1150# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X2955 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2956 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2957 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2958 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2959 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2960 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2961 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2962 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2964 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2965 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2966 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2967 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2968 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2970 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2971 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2972 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2973 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X2974 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2975 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2977 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2978 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2979 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2980 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2981 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2982 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2983 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2984 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2985 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2986 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X2987 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2988 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2989 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2990 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X2992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2994 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2995 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2996 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X2997 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2998 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X2999 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3000 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3001 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3003 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3004 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3005 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3007 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3008 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3009 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3010 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3011 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3012 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3013 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3014 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3015 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3016 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3017 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3018 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3020 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3021 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3022 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3023 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3024 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3026 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3027 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3028 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3030 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3031 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3032 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3034 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3035 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3036 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3037 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3038 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3039 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3040 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3041 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3042 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3044 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3045 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3046 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3047 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3048 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3049 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3050 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=5.5934 pd=16.02 as=2.0274 ps=14.09 w=4.38 l=0.5
X3051 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3052 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3053 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3054 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3055 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3056 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3057 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3058 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3059 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3060 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3061 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3062 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3063 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3064 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3065 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3066 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3067 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3068 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3069 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3070 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3071 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3072 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3073 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3074 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3075 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3076 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3077 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3078 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3079 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3081 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3082 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3083 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3084 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3085 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3086 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3087 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3088 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3089 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3090 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3091 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3093 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3095 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3096 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3097 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3098 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3100 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3101 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3103 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3104 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3105 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3106 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3107 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3109 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3111 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3112 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3113 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3114 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3115 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3116 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3117 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3118 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3119 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3120 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3121 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3122 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3123 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3125 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3126 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3127 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3128 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3129 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3130 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3131 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3132 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3133 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3134 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3135 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3137 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3138 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3139 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3140 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3141 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3142 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3143 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3144 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3147 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3148 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3149 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3150 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3153 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3154 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3155 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3156 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3157 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3158 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3159 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3163 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3165 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3166 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3167 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3168 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3169 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3170 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3173 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3174 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3175 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3176 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3177 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3178 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3179 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3180 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3181 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3182 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3185 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3186 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3187 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3189 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3190 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3191 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3192 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3193 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3194 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3195 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3196 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3198 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3199 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3200 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3201 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3202 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3203 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3205 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3207 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3208 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3209 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3210 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3211 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3212 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3214 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3215 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3216 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3217 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3218 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3219 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3221 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3222 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3224 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3226 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3227 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3228 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3229 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3230 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3231 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3232 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3233 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3234 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3235 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3236 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3237 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3238 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3239 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3240 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3241 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3243 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3244 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3246 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3247 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3248 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3249 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3250 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3251 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3252 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3254 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3255 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3256 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3257 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3259 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3260 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3262 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3263 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3265 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3266 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3267 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3269 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3270 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3271 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3274 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3275 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3276 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3278 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3279 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3284 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3286 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3288 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3289 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3290 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3291 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3292 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3293 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3294 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3295 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3296 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3298 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3299 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3300 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3301 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3303 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3306 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3307 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3308 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3309 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3310 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3311 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3312 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3314 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3315 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3316 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3317 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3320 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3321 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3324 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3325 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3326 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3327 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3328 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3329 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3330 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3332 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3333 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3334 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3335 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3336 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3337 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3339 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3340 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3341 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3342 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3343 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3344 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3345 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3347 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3348 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3349 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3350 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3351 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3352 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3353 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3354 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3355 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3356 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3360 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3361 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3362 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3363 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3364 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3365 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3367 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3368 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3369 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3370 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3371 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3373 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3374 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3375 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3376 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3377 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3378 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3379 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3380 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3381 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3382 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3383 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3384 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3385 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3386 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3387 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3389 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3393 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3394 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3395 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3396 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3397 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3400 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3401 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3402 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3403 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3404 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3405 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3406 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3408 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3410 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3411 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3412 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3413 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3414 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3415 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3417 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3419 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3420 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3421 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3422 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3424 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3425 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3426 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3427 a_112_1150# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X3428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3429 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3431 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3432 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3434 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3436 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3437 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3438 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3439 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3440 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3441 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3442 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3443 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3444 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3445 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3446 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3447 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3448 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3451 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3452 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3453 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3454 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3455 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3457 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3458 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3459 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3460 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3461 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3462 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3463 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3466 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3467 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3468 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3470 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3471 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3474 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3476 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3477 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3478 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3479 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3480 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3481 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3482 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3483 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3484 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3485 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3486 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3487 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3488 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3489 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3490 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3492 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3493 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3494 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3495 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3496 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3499 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3503 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3504 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3505 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3506 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3507 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3508 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3509 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3510 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3511 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3512 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3513 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3514 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3515 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3516 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3517 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3518 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3519 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3520 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3521 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3522 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3523 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3524 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3525 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3526 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3527 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3528 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3529 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3530 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3531 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3532 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3533 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3534 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3535 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3536 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3537 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3538 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3539 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3540 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3541 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3542 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3543 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3544 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3545 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3546 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3547 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3548 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3549 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3550 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3551 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3552 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3553 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3554 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3555 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3556 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3557 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3558 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3559 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3560 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3561 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3562 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3563 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3564 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3565 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3566 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3567 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3568 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3569 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3570 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3571 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3572 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3573 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3574 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3575 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3576 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3577 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3578 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3579 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3580 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3581 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3582 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3583 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3584 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3585 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3586 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3587 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3588 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3589 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3590 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3591 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3592 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3593 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3594 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3595 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3596 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3597 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3598 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3599 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3600 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3601 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3602 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3603 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3604 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3605 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3606 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3607 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3608 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3609 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3610 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3611 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3612 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3613 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3614 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3615 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3616 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3617 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3618 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3619 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3620 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3621 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3622 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3623 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3624 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3625 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3626 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3627 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3628 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3629 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3630 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3631 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3632 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3633 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3634 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3635 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3636 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3637 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3638 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3639 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3640 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3641 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3642 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3643 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3644 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3645 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3646 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3647 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3648 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3649 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3650 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3651 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3652 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3653 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3654 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3655 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3656 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3657 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3658 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3659 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3660 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3661 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3662 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3663 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3664 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3665 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3666 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3667 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3668 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3669 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3670 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3671 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3672 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3673 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3674 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3675 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3676 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3677 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3678 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3679 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3680 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3681 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3682 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3683 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3684 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3685 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3686 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3687 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3688 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3689 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3690 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3691 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3692 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3693 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3694 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3695 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3696 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3697 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3698 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3699 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3700 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3701 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3702 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3703 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3704 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3705 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3706 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3707 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3708 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3709 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3710 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3711 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3712 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3713 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3714 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3715 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3716 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3717 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3718 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3719 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3720 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3721 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3722 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3723 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3724 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3725 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3726 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3727 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3728 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3729 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3730 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3731 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3732 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3733 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3734 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3735 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3736 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3737 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3738 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3739 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3740 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3741 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3742 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3743 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3744 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3745 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3746 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3747 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3748 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3749 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3750 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3751 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3752 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3753 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3754 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3755 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3756 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3757 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3758 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3759 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3760 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3761 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3762 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3763 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3764 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3765 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3766 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3767 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3768 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3769 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3770 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3771 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3772 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3773 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3774 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3775 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3776 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3777 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3778 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3779 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3780 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3781 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3782 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3783 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3784 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3785 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3786 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3787 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3788 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3789 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3790 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3791 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3792 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3793 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3794 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3795 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3796 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3797 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3798 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3799 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3800 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3801 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3802 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3803 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3804 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3805 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3806 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3807 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3808 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3809 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3810 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3811 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3812 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3813 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3814 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3815 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3816 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3817 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3818 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3819 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3820 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3821 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3822 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3823 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3824 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3825 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3826 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3827 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3828 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3829 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3830 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3831 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3832 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3833 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3834 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3835 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3836 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3837 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3838 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3839 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3840 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3841 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3842 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3843 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3844 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3845 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3846 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3847 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3848 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3849 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3850 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3851 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3852 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3853 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3854 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3855 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3856 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3857 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3858 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3859 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3860 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3861 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3862 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3863 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3864 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3865 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3866 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3867 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3868 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3869 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3870 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3871 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3872 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3873 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3874 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3875 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3876 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3877 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3878 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3879 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3880 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3881 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3882 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3883 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3884 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3885 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3886 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3887 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3888 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3889 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3890 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3891 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3892 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3893 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3894 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3895 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3896 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3897 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3898 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3899 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3900 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3901 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3902 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3903 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3904 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3905 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X3906 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3907 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3908 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3909 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3910 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3911 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3912 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3913 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3914 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3915 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3916 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3917 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3918 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3919 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3920 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3921 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3922 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3923 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3924 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3925 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3926 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3927 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3928 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3929 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3930 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3931 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3932 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3933 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3934 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3935 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3936 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3937 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3938 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3939 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3940 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3941 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3942 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3943 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3944 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3945 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3946 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3947 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3948 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3949 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3950 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3951 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3952 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3953 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3954 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3955 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3956 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3957 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3958 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3959 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3960 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3961 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3962 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3963 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3964 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3965 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3966 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3967 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3968 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3969 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3970 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3971 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3972 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3973 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3974 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3975 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3976 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X3977 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3978 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3979 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3980 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3981 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3982 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X3983 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3984 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3985 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X3986 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3987 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3988 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3989 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3990 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3991 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3992 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3993 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X3994 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3995 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X3996 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3997 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X3998 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X3999 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4000 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4001 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4002 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4003 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4004 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4005 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4006 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4007 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4008 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4009 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4010 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4011 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4012 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4013 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4014 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4015 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4016 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4017 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4018 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4019 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4020 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4021 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4022 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4023 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4024 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4025 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4026 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4027 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4028 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4029 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4030 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4031 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4032 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4033 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4034 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4035 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4036 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4037 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4038 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4039 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4040 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4041 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4042 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4043 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4044 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4045 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4046 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4047 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4048 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4049 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4050 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4051 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4052 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4053 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4054 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4055 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4056 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4057 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4058 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4059 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4060 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4061 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4062 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4063 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4064 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4065 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4066 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4067 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4068 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4069 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4070 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4071 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4072 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4073 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4074 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4075 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4076 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4077 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4078 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4079 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4080 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4081 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4082 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4083 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4084 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4085 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4086 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4087 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4088 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4089 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4090 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4091 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4092 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4093 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4094 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4095 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4096 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4097 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4098 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4099 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4100 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4101 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4102 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4103 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4104 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4105 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4106 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4107 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4108 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4109 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4110 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4111 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4112 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4113 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4114 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4115 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4116 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4117 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4118 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4119 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4120 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4121 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4122 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4123 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4124 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4125 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4126 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4127 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4128 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4129 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4130 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4131 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4132 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4133 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4134 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4135 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4136 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4137 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4138 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4139 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4140 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4141 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4142 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4143 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4144 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4145 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4146 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4147 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4148 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4149 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4150 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4151 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4152 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4153 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4154 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4155 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.7846 ps=18.84 w=4.38 l=0.5
X4156 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4157 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4158 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4159 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4160 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4161 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4162 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4163 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4164 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4165 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4166 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4167 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4168 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4169 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4170 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4171 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4172 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4173 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4174 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4175 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4176 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4177 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4178 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4179 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4180 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4181 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4182 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4183 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4184 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4185 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4186 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4187 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4188 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4189 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4190 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4191 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4192 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4193 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4194 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4195 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4196 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4197 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4198 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4199 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4200 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4201 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4202 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4203 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4204 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4205 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4206 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4207 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4208 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4209 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4210 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4211 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4212 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4213 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4214 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4215 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4216 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4217 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4218 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4219 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4220 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4221 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4222 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4223 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4224 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4225 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4226 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4227 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4228 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4229 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4230 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4231 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4232 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4233 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4234 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4235 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4236 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4237 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4238 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4239 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4240 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4241 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4242 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4243 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4244 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4245 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4246 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4247 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4248 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4249 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4250 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4251 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4252 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4253 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4254 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4255 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4256 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4257 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4258 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4259 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4260 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4261 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4262 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4263 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4264 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4265 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4266 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4267 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4268 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4269 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4270 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4271 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4272 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4273 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4274 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4275 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4276 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4277 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4278 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4279 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4280 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4281 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4282 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4283 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4284 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4285 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4286 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4287 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4288 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4289 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4290 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4291 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4292 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4293 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4294 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4295 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4296 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4297 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4298 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4299 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4300 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4301 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4302 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4303 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4304 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4305 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4306 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4307 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4308 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4309 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4310 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4311 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4312 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4313 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4314 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4315 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4316 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4317 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4318 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4319 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4320 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4321 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4322 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4323 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4324 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4325 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4326 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4327 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4328 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4329 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4330 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4331 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4332 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4333 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4334 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4335 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4336 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4337 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4338 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4339 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4340 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4341 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4342 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4343 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4344 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4345 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4346 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4347 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4348 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4349 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4350 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4351 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4352 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4353 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4354 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4355 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4356 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4357 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4358 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4359 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4360 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4361 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4362 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4363 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4364 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4365 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4366 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4367 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4368 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4369 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4370 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4371 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4372 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4373 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4374 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4375 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4376 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4377 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4378 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4379 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4380 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4381 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4382 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4383 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4384 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4385 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4386 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4387 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4388 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4389 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4390 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4391 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4392 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4393 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4394 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4395 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4396 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4397 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4398 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4399 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4400 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4401 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4402 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4403 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4404 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4405 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4406 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4407 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4408 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4409 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4410 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4411 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4412 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.2285 ps=16.31 w=4.38 l=0.5
X4413 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4414 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4415 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4416 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4417 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4418 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4419 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4420 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4421 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4422 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4423 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4424 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4425 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4426 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4427 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4428 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4429 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4430 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4431 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4432 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4433 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4434 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4435 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4436 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4437 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4438 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4439 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4440 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4441 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4442 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4443 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4444 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4445 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4446 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4447 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4448 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4449 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4450 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4451 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4452 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4453 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4454 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4455 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4456 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4457 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4458 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4459 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4460 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4461 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4462 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4463 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4464 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4465 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4466 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4467 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4468 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4469 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4470 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4471 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4472 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4473 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4474 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4475 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4476 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4477 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4478 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4479 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4480 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4481 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4482 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.2285 pd=16.31 as=2.0274 ps=14.09 w=4.38 l=0.5
X4483 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4484 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4485 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.2285 ps=16.31 w=4.38 l=0.5
X4486 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4487 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4488 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4489 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4490 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4491 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4492 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4493 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.0274 ps=14.09 w=4.38 l=0.5
X4494 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4495 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4496 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4497 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4498 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4499 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4500 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4501 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4502 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4503 a_112_1150# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=5.5934 ps=16.02 w=4.38 l=0.5
X4504 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4505 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4506 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4507 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.0274 pd=14.09 as=6.8636 ps=16.6 w=4.38 l=0.5
X4508 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4509 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
X4510 dw_n11050_n11060# a_n50_n50# a_112_3350# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=6.8636 pd=16.6 as=2.7846 ps=18.84 w=4.38 l=0.5
X4511 a_112_3350# a_n50_n50# dw_n11050_n11060# dw_n11050_n11060# sky130_fd_pr__pfet_g5v0d10v5 ad=2.7846 pd=18.84 as=6.8636 ps=16.6 w=4.38 l=0.5
.ends

.subckt power_stage p_in sw_node vdd_pwr sky130_fd_sc_hd__inv_4_1/VPB vss dvss
Xsky130_fd_sc_hd__decap_3_0 dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_1 dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__inv_4_0 p_in dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ gate_drive_0/in_m sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_1 gate_drive_0/in_m dvss dvss sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__inv_4_1/VPB gate_drive_0/in_p sky130_fd_sc_hd__inv_4
Xgate_drive_0 gate_drive_0/in_m gate_drive_0/in_p gate_drive_0/out vdd_pwr vss dvss
+ gate_drive
Xsky130_fd_sc_hd__diode_2_0 p_in dvss dvss sky130_fd_sc_hd__inv_4_1/VPB sky130_fd_sc_hd__inv_4_1/VPB
+ sky130_fd_sc_hd__diode_2
Xpmos_waffle_48x48_0 vdd_pwr vss gate_drive_0/out sw_node sw_node pmos_waffle_48x48
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.178875 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.178875 ps=1.26 w=0.75 l=0.5
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ a_n3678_n531# a_296_n557# a_950_n531#
+ a_n2374_n557# a_3976_n531# a_2908_n531# a_n1306_n557# a_n3442_n557# a_n2076_n531#
+ a_n3144_n531# a_2610_n557# a_1542_n557# a_n950_n557# a_n1008_n531# a_n4212_n531#
+ a_3442_n531# a_2374_n531# a_1306_n531# a_n652_n531# a_1898_n557# a_n3798_n557# a_2966_n557#
+ a_772_n531# a_118_n557# a_3798_n531# a_n1720_n531# a_n1128_n557# a_n2196_n557# a_n3264_n557#
+ a_1364_n557# a_3500_n557# a_2432_n557# a_n772_n557# a_2196_n531# a_n474_n531# a_n4034_n531#
+ a_3264_n531# a_1128_n531# a_830_n557# a_3856_n557# a_2788_n557# a_n1840_n557# a_594_n531#
+ a_n1542_n531# a_n2610_n531# a_n3086_n557# a_2254_n557# a_1186_n557# a_n594_n557#
+ a_n2018_n557# a_n4154_n557# a_1840_n531# a_3322_n557# a_3086_n531# a_n296_n531#
+ a_n1898_n531# a_n2966_n531# a_4154_n531# a_2018_n531# a_60_n531# a_652_n557# a_3678_n557#
+ a_n1662_n557# a_n2730_n557# a_n1364_n531# a_n60_n557# a_416_n531# a_n2432_n531#
+ a_1662_n531# a_n3500_n531# a_3144_n557# a_2076_n557# a_1008_n557# a_2730_n531# a_n416_n557#
+ a_n2788_n531# a_n3856_n531# a_474_n557# a_n118_n531# a_n1484_n557# a_n2552_n557#
+ a_n3620_n557# a_238_n531# a_n1186_n531# a_n2254_n531# a_1720_n557# a_n3322_n531#
+ a_n4346_n691# a_2552_n531# a_1484_n531# a_n830_n531# a_4034_n557# a_n3976_n557#
+ a_3620_n531# a_n238_n557# a_n2908_n557#
X0 a_n3856_n531# a_n3976_n557# a_n4034_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_2196_n531# a_2076_n557# a_2018_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n2610_n531# a_n2730_n557# a_n2788_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n2254_n531# a_n2374_n557# a_n2432_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n652_n531# a_n772_n557# a_n830_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_2018_n531# a_1898_n557# a_1840_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n1008_n531# a_n1128_n557# a_n1186_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_594_n531# a_474_n557# a_416_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_3264_n531# a_3144_n557# a_3086_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n3322_n531# a_n3442_n557# a_n3500_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_60_n531# a_n60_n557# a_n118_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_3086_n531# a_2966_n557# a_2908_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_1484_n531# a_1364_n557# a_1306_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_n1542_n531# a_n1662_n557# a_n1720_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_2552_n531# a_2432_n557# a_2374_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_n3678_n531# a_n3798_n557# a_n3856_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_950_n531# a_830_n557# a_772_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X17 a_3620_n531# a_3500_n557# a_3442_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X18 a_n2076_n531# a_n2196_n557# a_n2254_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X19 a_n830_n531# a_n950_n557# a_n1008_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X20 a_n474_n531# a_n594_n557# a_n652_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X21 a_1840_n531# a_1720_n557# a_1662_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X22 a_n3500_n531# a_n3620_n557# a_n3678_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X23 a_416_n531# a_296_n557# a_238_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X24 a_n3144_n531# a_n3264_n557# a_n3322_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X25 a_2908_n531# a_2788_n557# a_2730_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X26 a_n1898_n531# a_n2018_n557# a_n2076_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X27 a_4154_n531# a_4034_n557# a_3976_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X28 a_n296_n531# a_n416_n557# a_n474_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 a_1306_n531# a_1186_n557# a_1128_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X30 a_3976_n531# a_3856_n557# a_3798_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X31 a_n1720_n531# a_n1840_n557# a_n1898_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X32 a_n1364_n531# a_n1484_n557# a_n1542_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X33 a_238_n531# a_118_n557# a_60_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X34 a_2374_n531# a_2254_n557# a_2196_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X35 a_n2788_n531# a_n2908_n557# a_n2966_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X36 a_n2432_n531# a_n2552_n557# a_n2610_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X37 a_1128_n531# a_1008_n557# a_950_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X38 a_n1186_n531# a_n1306_n557# a_n1364_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X39 a_772_n531# a_652_n557# a_594_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X40 a_3442_n531# a_3322_n557# a_3264_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 a_1662_n531# a_1542_n557# a_1484_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X42 a_n2966_n531# a_n3086_n557# a_n3144_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X43 a_2730_n531# a_2610_n557# a_2552_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X44 a_n4034_n531# a_n4154_n557# a_n4212_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X45 a_n118_n531# a_n238_n557# a_n296_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X46 a_3798_n531# a_3678_n557# a_3620_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY a_652_n562# a_n1186_n536# a_238_n536#
+ a_n1662_n562# a_3678_n562# a_n2254_n536# a_n2730_n562# a_n3322_n536# a_n60_n562#
+ a_1484_n536# a_2552_n536# a_n830_n536# a_3620_n536# w_n4412_n762# a_2076_n562# a_3144_n562#
+ a_1008_n562# a_n3678_n536# a_n416_n562# a_950_n536# a_474_n562# a_3976_n536# a_2908_n536#
+ a_n1484_n562# a_n2076_n536# a_n2552_n562# a_n3144_n536# a_n1008_n536# a_n3620_n562#
+ a_n4212_n536# a_1720_n562# a_2374_n536# a_n652_n536# a_1306_n536# a_3442_n536# a_n3976_n562#
+ a_4034_n562# a_n238_n562# a_772_n536# a_n2908_n562# a_296_n562# a_3798_n536# a_n1720_n536#
+ a_n2374_n562# a_n3442_n562# a_n1306_n562# a_n4034_n536# a_1542_n562# a_2196_n536#
+ a_n474_n536# a_2610_n562# a_n950_n562# a_1128_n536# a_3264_n536# a_n3798_n562# a_594_n536#
+ a_1898_n562# a_2966_n562# a_n1542_n536# a_n2610_n536# a_118_n562# a_n2196_n562#
+ a_1840_n536# a_n3264_n562# a_n1128_n562# a_1364_n562# a_n1898_n536# a_n296_n536#
+ a_2432_n562# a_n2966_n536# a_n772_n562# a_3086_n536# a_3500_n562# a_2018_n536# a_4154_n536#
+ a_60_n536# a_830_n562# a_2788_n562# a_n1364_n536# a_416_n536# a_n1840_n562# a_3856_n562#
+ a_n2432_n536# a_n3500_n536# a_1662_n536# a_n3086_n562# a_2730_n536# a_n4154_n562#
+ a_n2018_n562# a_1186_n562# a_2254_n562# a_n2788_n536# a_n594_n562# a_3322_n562#
+ a_n3856_n536# a_n118_n536#
X0 a_2552_n536# a_2432_n562# a_2374_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_950_n536# a_830_n562# a_772_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_3620_n536# a_3500_n562# a_3442_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n3678_n536# a_n3798_n562# a_n3856_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n830_n536# a_n950_n562# a_n1008_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n2076_n536# a_n2196_n562# a_n2254_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n474_n536# a_n594_n562# a_n652_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_1840_n536# a_1720_n562# a_1662_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_416_n536# a_296_n562# a_238_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n3500_n536# a_n3620_n562# a_n3678_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_n3144_n536# a_n3264_n562# a_n3322_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_2908_n536# a_2788_n562# a_2730_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_4154_n536# a_4034_n562# a_3976_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X13 a_n1898_n536# a_n2018_n562# a_n2076_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_n296_n536# a_n416_n562# a_n474_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_1306_n536# a_1186_n562# a_1128_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_n1720_n536# a_n1840_n562# a_n1898_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X17 a_n1364_n536# a_n1484_n562# a_n1542_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X18 a_238_n536# a_118_n562# a_60_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X19 a_3976_n536# a_3856_n562# a_3798_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X20 a_n2788_n536# a_n2908_n562# a_n2966_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X21 a_2374_n536# a_2254_n562# a_2196_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X22 a_n2432_n536# a_n2552_n562# a_n2610_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X23 a_1128_n536# a_1008_n562# a_950_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X24 a_n1186_n536# a_n1306_n562# a_n1364_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X25 a_772_n536# a_652_n562# a_594_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X26 a_3442_n536# a_3322_n562# a_3264_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X27 a_1662_n536# a_1542_n562# a_1484_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X28 a_n2966_n536# a_n3086_n562# a_n3144_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 a_2730_n536# a_2610_n562# a_2552_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X30 a_n4034_n536# a_n4154_n562# a_n4212_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X31 a_n118_n536# a_n238_n562# a_n296_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X32 a_3798_n536# a_3678_n562# a_3620_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X33 a_n3856_n536# a_n3976_n562# a_n4034_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X34 a_n2610_n536# a_n2730_n562# a_n2788_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X35 a_2196_n536# a_2076_n562# a_2018_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X36 a_n2254_n536# a_n2374_n562# a_n2432_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X37 a_n652_n536# a_n772_n562# a_n830_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X38 a_2018_n536# a_1898_n562# a_1840_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X39 a_n1008_n536# a_n1128_n562# a_n1186_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X40 a_594_n536# a_474_n562# a_416_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 a_3264_n536# a_3144_n562# a_3086_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X42 a_n3322_n536# a_n3442_n562# a_n3500_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X43 a_60_n536# a_n60_n562# a_n118_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X44 a_3086_n536# a_2966_n562# a_2908_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X45 a_1484_n536# a_1364_n562# a_1306_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X46 a_n1542_n536# a_n1662_n562# a_n1720_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ a_n919_n536# a_207_n562# a_n1217_n562#
+ w_n1653_n762# a_n385_n536# a_1039_n536# a_n861_n562# a_n1453_n536# a_505_n536# a_1275_n562#
+ a_29_n562# a_n1039_n562# a_n683_n562# a_n207_n536# a_741_n562# a_327_n536# a_n1275_n536#
+ a_1097_n562# a_n505_n562# a_n29_n536# a_n1097_n536# a_563_n562# a_149_n536# a_1395_n536#
+ a_n741_n536# a_919_n562# a_861_n536# a_n327_n562# a_385_n562# a_n1395_n562# a_1217_n536#
+ a_n563_n536# a_683_n536# a_n149_n562#
X0 a_n207_n536# a_n327_n562# a_n385_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_1217_n536# a_1097_n562# a_1039_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n1275_n536# a_n1395_n562# a_n1453_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X3 a_n741_n536# a_n861_n562# a_n919_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n1097_n536# a_n1217_n562# a_n1275_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_683_n536# a_563_n562# a_505_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_1039_n536# a_919_n562# a_861_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_n29_n536# a_n149_n562# a_n207_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n563_n536# a_n683_n562# a_n741_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n919_n536# a_n1039_n562# a_n1097_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_505_n536# a_385_n562# a_327_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_n385_n536# a_n505_n562# a_n563_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_1395_n536# a_1275_n562# a_1217_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X13 a_327_n536# a_207_n562# a_149_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_149_n536# a_29_n562# a_n29_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_861_n536# a_741_n562# a_683_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_CZUCEE a_4017_n2176# a_n9969_1744# a_8553_1744#
+ a_n6567_1744# a_n17151_1744# a_5151_1744# a_n3165_1744# a_16869_1744# a_13467_1744#
+ a_10065_1744# a_19137_n2176# a_17247_1744# a_2127_n2176# a_237_1744# a_n519_1744#
+ a_19515_n2176# a_n16017_n2176# a_2505_n2176# a_n9213_n2176# a_17247_n2176# a_n10725_1744#
+ a_n5811_1744# a_n9591_1744# a_n17907_1744# a_8175_n2176# a_9687_1744# a_5907_1744#
+ a_n14505_1744# a_n18285_1744# a_17625_n2176# a_6285_1744# a_2505_1744# a_n11103_1744#
+ a_n14127_n2176# a_12711_1744# a_16491_1744# a_n4299_1744# a_n7323_n2176# a_15357_n2176#
+ a_8553_n2176# a_11199_1744# a_n5055_n2176# a_n7701_n2176# a_n8079_1744# a_n14505_n2176#
+ a_13089_n2176# a_15735_n2176# a_6285_n2176# a_n141_n2176# a_n519_n2176# a_n141_1744#
+ a_n5433_n2176# a_n12237_n2176# a_8931_n2176# a_13467_n2176# a_6663_n2176# a_n3165_n2176#
+ a_n12615_n2176# a_11199_n2176# a_n5811_n2176# a_n11859_1744# a_n19927_n2306# a_13845_n2176#
+ a_4395_n2176# a_8931_1744# a_n3543_n2176# a_n10347_n2176# a_n6945_1744# a_n3543_1744#
+ a_n15639_1744# a_11577_n2176# a_3639_1744# a_n12237_1744# a_n18285_n2176# a_13845_1744#
+ a_4773_n2176# a_n1275_n2176# a_10443_1744# a_n10725_n2176# a_n897_1744# a_n3921_n2176#
+ a_n7323_1744# a_n19419_1744# a_11955_n2176# a_7419_1744# a_615_1744# a_n16017_1744#
+ a_17625_1744# a_4017_1744# a_n1653_n2176# a_n18663_n2176# a_14223_1744# a_n9591_n2176#
+ a_n16395_n2176# a_2883_n2176# a_n9969_n2176# a_18003_1744# a_2883_1744# a_n14883_1744#
+ a_n11481_1744# a_n16773_n2176# a_18003_n2176# a_n18663_1744# a_6663_1744# a_n4677_1744#
+ a_n15261_1744# a_3261_1744# a_n1275_1744# a_9309_n2176# a_14979_1744# a_11577_1744#
+ a_n14883_n2176# a_n19041_1744# a_16113_n2176# a_7041_1744# a_n897_n2176# a_n8457_1744#
+ a_n5055_1744# a_18759_1744# a_15357_1744# a_7419_n2176# a_7041_n2176# a_237_n2176#
+ a_n12993_n2176# a_19137_1744# a_14223_n2176# a_615_n2176# a_n3921_1744# a_14601_n2176#
+ a_5529_n2176# a_5151_n2176# a_n12615_1744# a_n19797_1744# a_7797_1744# a_993_1744#
+ a_n11103_n2176# a_n16395_1744# a_10821_1744# a_4395_1744# a_12333_n2176# a_n7701_1744#
+ a_n19041_n2176# a_n19419_n2176# a_5907_n2176# a_n2031_n2176# a_n2409_n2176# a_8175_1744#
+ a_10065_n2176# a_14601_1744# a_n2409_1744# a_n6189_1744# a_18381_1744# a_3261_n2176#
+ a_12711_n2176# a_3639_n2176# a_13089_1744# a_10443_n2176# a_n8079_n2176# a_n17151_n2176#
+ a_n17529_n2176# a_18381_n2176# a_18759_n2176# a_1749_n2176# a_1371_n2176# a_n8457_n2176#
+ a_10821_n2176# a_n17907_n2176# a_n6189_n2176# a_9687_n2176# a_n1653_1744# a_n13749_1744#
+ a_1749_1744# a_n8835_n2176# a_n10347_1744# a_n15261_n2176# a_n15639_n2176# a_11955_1744#
+ a_16491_n2176# a_16869_n2176# a_n8835_1744# a_n5433_1744# a_n6567_n2176# a_5529_1744#
+ a_n2031_1744# a_n17529_1744# a_15735_1744# a_2127_1744# a_n14127_1744# a_12333_1744#
+ a_n4299_n2176# a_7797_n2176# a_n6945_n2176# a_n13371_n2176# a_n13749_n2176# a_n9213_1744#
+ a_9309_1744# a_14979_n2176# a_19515_1744# a_993_n2176# a_16113_1744# a_n4677_n2176#
+ a_n12993_1744# a_n11481_n2176# a_n11859_n2176# a_n16773_1744# a_4773_1744# a_n13371_1744#
+ a_1371_1744# a_n2787_1744# a_n2787_n2176# a_n19797_n2176#
X0 a_n19419_1744# a_n19419_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X1 a_n19041_1744# a_n19041_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X2 a_993_1744# a_993_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X3 a_n16017_1744# a_n16017_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X4 a_9687_1744# a_9687_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X5 a_6285_1744# a_6285_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X6 a_18759_1744# a_18759_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X7 a_8553_1744# a_8553_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X8 a_5529_1744# a_5529_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X9 a_13089_1744# a_13089_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X10 a_n16773_1744# a_n16773_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X11 a_18381_1744# a_18381_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X12 a_n13749_1744# a_n13749_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X13 a_15357_1744# a_15357_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X14 a_5151_1744# a_5151_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X15 a_2127_1744# a_2127_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X16 a_17625_1744# a_17625_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X17 a_n9969_1744# a_n9969_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X18 a_n4299_1744# a_n4299_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X19 a_n10347_1744# a_n10347_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X20 a_n13371_1744# a_n13371_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X21 a_n6567_1744# a_n6567_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X22 a_n9591_1744# a_n9591_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X23 a_n12615_1744# a_n12615_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X24 a_14223_1744# a_14223_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X25 a_n8835_1744# a_n8835_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X26 a_n3165_1744# a_n3165_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X27 a_n5433_1744# a_n5433_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X28 a_n897_1744# a_n897_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X29 a_n2409_1744# a_n2409_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X30 a_n7701_1744# a_n7701_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X31 a_2883_1744# a_2883_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X32 a_n2031_1744# a_n2031_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X33 a_11955_1744# a_11955_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X34 a_10821_1744# a_10821_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X35 a_n19797_1744# a_n19797_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X36 a_8175_1744# a_8175_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X37 a_7419_1744# a_7419_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X38 a_n16395_1744# a_n16395_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X39 a_n18663_1744# a_n18663_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X40 a_n15639_1744# a_n15639_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X41 a_n17907_1744# a_n17907_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X42 a_17247_1744# a_17247_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X43 a_7041_1744# a_7041_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X44 a_4017_1744# a_4017_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X45 a_19515_1744# a_19515_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X46 a_n6189_1744# a_n6189_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X47 a_n12237_1744# a_n12237_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X48 a_n15261_1744# a_n15261_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X49 a_n8457_1744# a_n8457_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X50 a_n14505_1744# a_n14505_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X51 a_16113_1744# a_16113_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X52 a_n5055_1744# a_n5055_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X53 a_n11103_1744# a_n11103_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X54 a_n7323_1744# a_n7323_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X55 a_14979_1744# a_14979_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X56 a_4773_1744# a_4773_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X57 a_1749_1744# a_1749_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X58 a_n12993_1744# a_n12993_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X59 a_11577_1744# a_11577_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X60 a_1371_1744# a_1371_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X61 a_13845_1744# a_13845_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X62 a_n2787_1744# a_n2787_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X63 a_10443_1744# a_10443_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X64 a_12711_1744# a_12711_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X65 a_n1653_1744# a_n1653_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X66 a_615_1744# a_615_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X67 a_n3921_1744# a_n3921_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X68 a_9309_1744# a_9309_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X69 a_n18285_1744# a_n18285_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X70 a_n17529_1744# a_n17529_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X71 a_19137_1744# a_19137_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X72 a_n17151_1744# a_n17151_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X73 a_n8079_1744# a_n8079_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X74 a_n14127_1744# a_n14127_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X75 a_18003_1744# a_18003_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X76 a_7797_1744# a_7797_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X77 a_n9213_1744# a_n9213_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X78 a_4395_1744# a_4395_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X79 a_16869_1744# a_16869_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X80 a_6663_1744# a_6663_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X81 a_3639_1744# a_3639_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X82 a_11199_1744# a_11199_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X83 a_8931_1744# a_8931_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X84 a_5907_1744# a_5907_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X85 a_n519_1744# a_n519_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X86 a_16491_1744# a_16491_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X87 a_n11859_1744# a_n11859_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X88 a_n14883_1744# a_n14883_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X89 a_13467_1744# a_13467_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X90 a_3261_1744# a_3261_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X91 a_15735_1744# a_15735_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X92 a_2505_1744# a_2505_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X93 a_n141_1744# a_n141_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X94 a_10065_1744# a_10065_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X95 a_n11481_1744# a_n11481_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X96 a_n4677_1744# a_n4677_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X97 a_n10725_1744# a_n10725_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X98 a_12333_1744# a_12333_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X99 a_14601_1744# a_14601_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X100 a_n6945_1744# a_n6945_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X101 a_n1275_1744# a_n1275_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X102 a_n3543_1744# a_n3543_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X103 a_237_1744# a_237_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
X104 a_n5811_1744# a_n5811_n2176# a_n19927_n2306# sky130_fd_pr__res_xhigh_po_1p41 l=17.6
.ends

.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
.ends

.subckt rstring_mux_ov vout ena otrip_decoded_avdd[15] otrip_decoded_avdd[14] otrip_decoded_avdd[13]
+ otrip_decoded_avdd[12] otrip_decoded_avdd[11] otrip_decoded_avdd[10] otrip_decoded_avdd[9]
+ otrip_decoded_avdd[8] otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5]
+ otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1]
+ otrip_decoded_avdd[0] vtop avdd avss
Xsky130_fd_pr__nfet_g5v0d10v5_K8JYEQ_0 vout otrip_decoded_avdd[8] vout otrip_decoded_avdd[3]
+ vtrip15 vtrip13 otrip_decoded_avdd[5] otrip_decoded_avdd[1] vout vout avss avss
+ otrip_decoded_avdd[6] vout vout vtrip14 vtrip12 vtrip10 vout otrip_decoded_avdd[11]
+ avss otrip_decoded_avdd[13] vtrip9 otrip_decoded_avdd[8] vout vout avss avss avss
+ otrip_decoded_avdd[10] otrip_decoded_avdd[14] otrip_decoded_avdd[12] otrip_decoded_avdd[6]
+ vout vout vtrip0 vout vout otrip_decoded_avdd[9] otrip_decoded_avdd[15] otrip_decoded_avdd[13]
+ otrip_decoded_avdd[4] vout vout vout otrip_decoded_avdd[2] otrip_decoded_avdd[12]
+ otrip_decoded_avdd[10] avss otrip_decoded_avdd[4] otrip_decoded_avdd[0] vtrip11
+ otrip_decoded_avdd[14] vout vtrip7 vtrip4 vtrip2 vout vout vout otrip_decoded_avdd[9]
+ avss avss avss vtrip5 avss vout vtrip3 vout vtrip1 avss avss avss vout otrip_decoded_avdd[7]
+ vout vout avss vout otrip_decoded_avdd[5] otrip_decoded_avdd[3] otrip_decoded_avdd[1]
+ vtrip8 vout vout otrip_decoded_avdd[11] vout avss vout vout vtrip6 otrip_decoded_avdd[15]
+ otrip_decoded_avdd[0] vout otrip_decoded_avdd[7] otrip_decoded_avdd[2] sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ
Xsky130_fd_pr__pfet_g5v0d10v5_4Z8MHY_0 otrip_decoded_b_avdd[9] vout vtrip8 avdd avdd
+ vout avdd vout avdd vout vout vtrip6 vout avdd avdd avdd avdd vout otrip_decoded_b_avdd[7]
+ vout avdd vtrip15 vtrip13 otrip_decoded_b_avdd[5] vout otrip_decoded_b_avdd[3] vout
+ vout otrip_decoded_b_avdd[1] vout otrip_decoded_b_avdd[11] vtrip12 vout vtrip10
+ vtrip14 otrip_decoded_b_avdd[0] sky130_fd_sc_hvl__inv_1_0[15]/Y otrip_decoded_b_avdd[7]
+ vtrip9 otrip_decoded_b_avdd[2] otrip_decoded_b_avdd[8] vout vout otrip_decoded_b_avdd[3]
+ otrip_decoded_b_avdd[1] otrip_decoded_b_avdd[5] vtrip0 avdd vout vout avdd otrip_decoded_b_avdd[6]
+ vout vout avdd vout otrip_decoded_b_avdd[11] otrip_decoded_b_avdd[13] vout vout
+ otrip_decoded_b_avdd[8] avdd vtrip11 avdd avdd otrip_decoded_b_avdd[10] vtrip4 vtrip7
+ otrip_decoded_b_avdd[12] vtrip2 otrip_decoded_b_avdd[6] vout otrip_decoded_b_avdd[14]
+ vout vout vout otrip_decoded_b_avdd[9] otrip_decoded_b_avdd[13] vtrip5 vout otrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1_0[15]/Y vtrip3 vtrip1 vout otrip_decoded_b_avdd[2] vout
+ otrip_decoded_b_avdd[0] otrip_decoded_b_avdd[4] otrip_decoded_b_avdd[10] otrip_decoded_b_avdd[12]
+ vout avdd otrip_decoded_b_avdd[14] vout vout sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY
Xsky130_fd_pr__pfet_g5v0d10v5_WY4TLZ_0 vtop ena_b ena_b avdd avdd avdd ena_b avdd
+ vtop ena_b ena_b ena_b ena_b vtop ena_b avdd vtop ena_b ena_b avdd avdd ena_b vtop
+ avdd avdd ena_b vtop ena_b ena_b ena_b vtop vtop avdd ena_b sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ
Xsky130_fd_pr__res_xhigh_po_1p41_CZUCEE_0 m1_12242_140# m1_n1744_4059# vtrip9 m1_2036_4059#
+ m1_n8548_4059# m1_13376_4059# m1_5060_4059# m1_25472_4059# m1_21692_4059# vtrip13
+ m1_27362_140# m1_25472_4059# m1_10730_140# m1_8840_4059# m1_8084_4059# avss m1_n7414_140#
+ m1_10730_140# m1_n610_140# m1_25850_140# m1_n2500_4059# m1_2792_4059# m1_n988_4059#
+ m1_n9304_4059# vtrip8 vtrip11 vtrip1 m1_n6280_4059# m1_n10060_4059# m1_25850_140#
+ vtrip3 m1_11108_4059# m1_n2500_4059# m1_n5902_140# m1_20936_4059# m1_24716_4059#
+ m1_4304_4059# m1_902_140# m1_23582_140# vtrip8 vtrip15 m1_3170_140# m1_902_140#
+ m1_524_4059# m1_n5902_140# m1_21314_140# m1_24338_140# vtrip2 m1_8462_140# m1_7706_140#
+ m1_8084_4059# m1_3170_140# m1_n3634_140# vtrip10 m1_22070_140# vtrip4 m1_5438_140#
+ m1_n4390_140# m1_19802_140# m1_2414_140# m1_n3256_4059# avss m1_22070_140# m1_12998_140#
+ vtrip9 m1_4682_140# m1_n2122_140# m1_1280_4059# m1_5060_4059# m1_n7036_4059# m1_19802_140#
+ m1_11864_4059# m1_n4012_4059# m1_n9682_140# m1_22448_4059# m1_12998_140# m1_6950_140#
+ vtrip13 m1_n2122_140# m1_7328_4059# m1_4682_140# m1_1280_4059# m1_n10816_4059# m1_20558_140#
+ vtrip5 m1_8840_4059# m1_n7792_4059# m1_26228_4059# m1_12620_4059# m1_6950_140# m1_n10438_140#
+ m1_22448_4059# m1_n1366_140# m1_n8170_140# m1_11486_140# m1_n1366_140# m1_26228_4059#
+ m1_11108_4059# m1_n6280_4059# m1_n3256_4059# m1_n8170_140# m1_26606_140# m1_n10060_4059#
+ vtrip3 m1_3548_4059# m1_n7036_4059# m1_11864_4059# m1_7328_4059# vtrip10 m1_23204_4059#
+ m1_20180_4059# m1_n6658_140# m1_n10816_4059# m1_24338_140# vtrip5 m1_7706_140# m1_n232_4059#
+ m1_3548_4059# m1_26984_4059# m1_23960_4059# vtrip6 vtrip4 m1_8462_140# m1_n4390_140#
+ m1_27740_4059# m1_22826_140# m1_9218_140# m1_4304_4059# m1_22826_140# vtrip0 vtrip0
+ m1_n4012_4059# vtop vtrip7 m1_9596_4059# m1_n2878_140# m1_n7792_4059# vtrip15 m1_12620_4059#
+ m1_20558_140# m1_524_4059# m1_n10438_140# m1_n11194_140# vtrip2 m1_6194_140# m1_6194_140#
+ vtrip7 vtrip12 m1_23204_4059# m1_5816_4059# m1_2036_4059# m1_26984_4059# m1_11486_140#
+ m1_21314_140# m1_12242_140# m1_21692_4059# vtrip14 m1_146_140# m1_n8926_140# m1_n8926_140#
+ m1_26606_140# m1_27362_140# m1_9974_140# m1_9974_140# m1_146_140# vtrip14 m1_n9682_140#
+ m1_2414_140# vtrip12 m1_6572_4059# m1_n5524_4059# m1_10352_4059# m1_n610_140# m1_n1744_4059#
+ m1_n6658_140# m1_n7414_140# m1_20180_4059# m1_25094_140# m1_25094_140# m1_n232_4059#
+ m1_2792_4059# m1_1658_140# vtrip1 m1_6572_4059# m1_n9304_4059# m1_23960_4059# m1_10352_4059#
+ m1_n5524_4059# m1_20936_4059# m1_3926_140# vtrip6 m1_1658_140# m1_n5146_140# m1_n5146_140#
+ m1_n988_4059# vtrip11 m1_23582_140# m1_27740_4059# m1_9218_140# m1_24716_4059# m1_3926_140#
+ m1_n4768_4059# m1_n2878_140# m1_n3634_140# m1_n8548_4059# m1_13376_4059# m1_n4768_4059#
+ m1_9596_4059# m1_5816_4059# m1_5438_140# m1_n11194_140# sky130_fd_pr__res_xhigh_po_1p41_CZUCEE
Xsky130_fd_sc_hvl__inv_1_0[0] otrip_decoded_avdd[0] avss avss avdd avdd otrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[1] otrip_decoded_avdd[1] avss avss avdd avdd otrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[2] otrip_decoded_avdd[2] avss avss avdd avdd otrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[3] otrip_decoded_avdd[3] avss avss avdd avdd otrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[4] otrip_decoded_avdd[4] avss avss avdd avdd otrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[5] otrip_decoded_avdd[5] avss avss avdd avdd otrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[6] otrip_decoded_avdd[6] avss avss avdd avdd otrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[7] otrip_decoded_avdd[7] avss avss avdd avdd otrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[8] otrip_decoded_avdd[8] avss avss avdd avdd otrip_decoded_b_avdd[8]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[9] otrip_decoded_avdd[9] avss avss avdd avdd otrip_decoded_b_avdd[9]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[10] otrip_decoded_avdd[10] avss avss avdd avdd otrip_decoded_b_avdd[10]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[11] otrip_decoded_avdd[11] avss avss avdd avdd otrip_decoded_b_avdd[11]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[12] otrip_decoded_avdd[12] avss avss avdd avdd otrip_decoded_b_avdd[12]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[13] otrip_decoded_avdd[13] avss avss avdd avdd otrip_decoded_b_avdd[13]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[14] otrip_decoded_avdd[14] avss avss avdd avdd otrip_decoded_b_avdd[14]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[15] otrip_decoded_avdd[15] avss avss avdd avdd sky130_fd_sc_hvl__inv_1_0[15]/Y
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_1 ena avss avss avdd avdd ena_b sky130_fd_sc_hvl__inv_1
Xsky130_fd_pr__nfet_g5v0d10v5_CD9S2Z_0 avss avss vtop ena_b sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XZ4X25 a_n887_n588# a_n429_n588# a_487_n588#
+ a_n945_n500# a_29_n588# a_n487_n500# a_n1079_n722# a_n29_n500# a_887_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_887_n500# a_487_n588# a_429_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X3 a_n487_n500# a_n887_n588# a_n945_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP a_n1174_n500# a_n200_n597# a_200_n500#
+ a_n1116_n597# a_n716_n500# a_n258_n500# w_n1374_n797# a_1116_n500# a_n658_n597#
+ a_658_n500# a_716_n597# a_258_n597#
X0 a_1116_n500# a_716_n597# a_658_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1 a_200_n500# a_n200_n597# a_n258_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_n716_n500# a_n1116_n597# a_n1174_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X3 a_658_n500# a_258_n597# a_200_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 a_n258_n500# a_n658_n597# a_n716_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_62W3XE a_358_n500# a_158_n588# a_100_n500# a_n158_n500#
+ a_n358_n588# a_n100_n588# a_n550_n722# a_n416_n500#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_n158_n500# a_n358_n588# a_n416_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X2 a_358_n500# a_158_n588# a_100_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EC8RE7 a_416_n500# a_n1364_n500# a_830_n588#
+ a_n1676_n722# a_n118_n500# a_1186_n588# a_n594_n588# a_238_n500# a_n1186_n500# a_652_n588#
+ a_1484_n500# a_n830_n500# a_n60_n588# a_950_n500# a_1008_n588# a_n416_n588# a_n1008_n500#
+ a_474_n588# a_n1484_n588# a_n652_n500# a_772_n500# a_n238_n588# a_296_n588# a_n474_n500#
+ a_1128_n500# a_n1306_n588# a_n950_n588# a_594_n500# a_n1542_n500# a_n296_n500# a_118_n588#
+ a_60_n500# a_1364_n588# a_n1128_n588# a_n772_n588#
X0 a_416_n500# a_296_n588# a_238_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_n296_n500# a_n416_n588# a_n474_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_1306_n500# a_1186_n588# a_1128_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n1364_n500# a_n1484_n588# a_n1542_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X4 a_238_n500# a_118_n588# a_60_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_1128_n500# a_1008_n588# a_950_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n1186_n500# a_n1306_n588# a_n1364_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_772_n500# a_652_n588# a_594_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n118_n500# a_n238_n588# a_n296_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n652_n500# a_n772_n588# a_n830_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_n1008_n500# a_n1128_n588# a_n1186_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_594_n500# a_474_n588# a_416_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_60_n500# a_n60_n588# a_n118_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_1484_n500# a_1364_n588# a_1306_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X14 a_950_n500# a_830_n588# a_772_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_n830_n500# a_n950_n588# a_n1008_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_n474_n500# a_n594_n588# a_n652_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_75AJMX a_n3403_n597# a_5977_n500# a_5177_n597#
+ a_29_n597# a_n2603_n500# a_5119_n500# a_3461_n597# a_3403_n500# a_n6035_n500# a_n2545_n597#
+ a_n1745_n500# a_4319_n597# a_2545_n500# a_2603_n597# a_n5177_n500# a_n1687_n597#
+ a_n4261_n597# a_n887_n500# w_n6235_n797# a_n3461_n500# a_n5977_n597# a_n29_n500#
+ a_n5119_n597# a_1687_n500# a_1745_n597# a_n829_n597# a_4261_n500# a_887_n597# a_829_n500#
+ a_n4319_n500#
X0 a_3403_n500# a_2603_n597# a_2545_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1 a_n29_n500# a_n829_n597# a_n887_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_n5177_n500# a_n5977_n597# a_n6035_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X3 a_2545_n500# a_1745_n597# a_1687_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_4261_n500# a_3461_n597# a_3403_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_n4319_n500# a_n5119_n597# a_n5177_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X6 a_829_n500# a_29_n597# a_n29_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X7 a_n2603_n500# a_n3403_n597# a_n3461_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X8 a_1687_n500# a_887_n597# a_829_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X9 a_5119_n500# a_4319_n597# a_4261_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X10 a_n3461_n500# a_n4261_n597# a_n4319_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X11 a_n1745_n500# a_n2545_n597# a_n2603_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X12 a_5977_n500# a_5177_n597# a_5119_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X13 a_n887_n500# a_n1687_n597# a_n1745_n500# w_n6235_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP a_n358_n597# a_358_n500# a_n100_n597#
+ a_100_n500# a_n158_n500# a_158_n597# w_n616_n797# a_n416_n500#
X0 a_358_n500# a_158_n597# a_100_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_100_n500# a_n100_n597# a_n158_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n158_n500# a_n358_n597# a_n416_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QZVU2P a_2974_n500# a_2116_n500# a_n458_n500#
+ a_n2974_n588# a_n3032_n500# a_n2116_n588# a_n400_n588# a_1258_n500# a_2174_n588#
+ a_n2174_n500# a_n3166_n722# a_n1258_n588# a_1316_n588# a_458_n588# a_400_n500# a_n1316_n500#
X0 a_n2174_n500# a_n2974_n588# a_n3032_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1 a_1258_n500# a_458_n588# a_400_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_n1316_n500# a_n2116_n588# a_n2174_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X3 a_n458_n500# a_n1258_n588# a_n1316_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_2116_n500# a_1316_n588# a_1258_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_2974_n500# a_2174_n588# a_2116_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X6 a_400_n500# a_n400_n588# a_n458_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DVQADA a_48_n3916# a_n330_n3916# a_n708_n3916#
+ a_1182_3484# a_n2598_3484# a_n3354_n3916# a_n1086_n3916# a_n3732_n3916# a_n1464_n3916#
+ a_2694_n3916# a_n1842_n3916# a_n3862_n4046# a_1938_3484# a_48_3484# a_n1842_3484#
+ a_n2220_3484# a_2316_3484# a_426_n3916# a_1560_3484# a_n2976_3484# a_804_n3916#
+ a_n3354_3484# a_3072_n3916# a_426_3484# a_n2220_n3916# a_3450_n3916# a_n708_3484#
+ a_2694_3484# a_1182_n3916# a_1938_n3916# a_1560_n3916# a_3072_3484# a_n1086_3484#
+ a_n330_3484# a_n2598_n3916# a_n3732_3484# a_804_3484# a_n2976_n3916# a_2316_n3916#
+ a_3450_3484# a_n1464_3484#
X0 a_n330_3484# a_n330_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 a_3072_3484# a_3072_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 a_2316_3484# a_2316_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X3 a_n1086_3484# a_n1086_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 a_n3354_3484# a_n3354_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 a_n2220_3484# a_n2220_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X6 a_1938_3484# a_1938_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X7 a_2694_3484# a_2694_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X8 a_1560_3484# a_1560_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X9 a_n2976_3484# a_n2976_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X10 a_48_3484# a_48_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X11 a_n1842_3484# a_n1842_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X12 a_804_3484# a_804_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X13 a_n708_3484# a_n708_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 a_1182_3484# a_1182_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 a_n2598_3484# a_n2598_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X16 a_3450_3484# a_3450_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X17 a_n3732_3484# a_n3732_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X18 a_n1464_3484# a_n1464_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X19 a_426_3484# a_426_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7JLQGA a_416_n500# a_n238_n597# a_n118_n500#
+ a_296_n597# a_238_n500# a_n830_n500# a_118_n597# a_n772_n597# w_n1030_n797# a_772_n500#
+ a_n474_n500# a_n594_n597# a_652_n597# a_n60_n597# a_n296_n500# a_60_n500# a_n416_n597#
+ a_474_n597#
X0 a_n474_n500# a_n594_n597# a_n652_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_416_n500# a_296_n597# a_238_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n296_n500# a_n416_n597# a_n474_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_238_n500# a_118_n597# a_60_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_772_n500# a_652_n597# a_594_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n118_n500# a_n238_n597# a_n296_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n652_n500# a_n772_n597# a_n830_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X7 a_594_n500# a_474_n597# a_416_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_60_n500# a_n60_n597# a_n118_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3DCHX4 a_n1687_n1687# a_n3287_n557# a_29_599#
+ a_1629_1781# a_1687_n2869# a_n3287_n1713# a_3287_n2843# a_3287_n531# a_n1629_1755#
+ a_1687_n1713# a_n1687_n531# a_n1687_625# a_29_n2869# a_n3345_n2843# a_n1687_n2843#
+ a_1687_1755# a_29_n1713# a_n29_n531# a_3287_1781# a_29_1755# a_n29_n1687# a_n3345_625#
+ a_n3479_n3003# a_n1687_1781# a_1629_n1687# a_n29_625# a_n3287_1755# a_n1629_n557#
+ a_3287_625# a_1687_599# a_n3345_n531# a_1629_n531# a_n3287_599# a_n1629_n2869# a_3287_n1687#
+ a_n29_1781# a_1629_625# a_n29_n2843# a_1687_n557# a_n1629_n1713# a_n1629_599# a_1629_n2843#
+ a_29_n557# a_n3287_n2869# a_n3345_n1687# a_n3345_1781#
X0 a_n1687_625# a_n3287_599# a_n3345_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X1 a_1629_n531# a_29_n557# a_n29_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X2 a_1629_1781# a_29_1755# a_n29_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X3 a_3287_n531# a_1687_n557# a_1629_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X4 a_3287_1781# a_1687_1755# a_1629_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X5 a_n1687_n531# a_n3287_n557# a_n3345_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X6 a_n29_625# a_n1629_599# a_n1687_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X7 a_n1687_n1687# a_n3287_n1713# a_n3345_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X8 a_n1687_1781# a_n3287_1755# a_n3345_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X9 a_1629_n1687# a_29_n1713# a_n29_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X10 a_n1687_n2843# a_n3287_n2869# a_n3345_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X11 a_3287_n1687# a_1687_n1713# a_1629_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X12 a_1629_n2843# a_29_n2869# a_n29_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X13 a_1629_625# a_29_599# a_n29_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X14 a_3287_625# a_1687_599# a_1629_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X15 a_n29_n531# a_n1629_n557# a_n1687_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X16 a_3287_n2843# a_1687_n2869# a_1629_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X17 a_n29_1781# a_n1629_1755# a_n1687_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X18 a_n29_n1687# a_n1629_n1713# a_n1687_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X19 a_n29_n2843# a_n1629_n2869# a_n1687_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
.ends

.subckt ibias_gen_ov itest ibias ibg_200n vbg_1v2 isrc_sel ena ve avss avdd
Xsky130_fd_pr__nfet_g5v0d10v5_XZ4X25_0 isrc_sel_b ena_b isrc_sel avss ena_b vn1 avss
+ avss avss vn0 sky130_fd_pr__nfet_g5v0d10v5_XZ4X25
Xsky130_fd_pr__pfet_g5v0d10v5_Y9S9FP_0 avdd ena vp0 isrc_sel vp1 avdd avdd vp ena
+ avdd ena isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP
Xsky130_fd_pr__nfet_g5v0d10v5_62W3XE_0 avss isrc_sel isrc_sel_b ena_b ena avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_62W3XE
Xsky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1 vp0 vstart isrc_sel avss vn0 isrc_sel vbg_1v2
+ vn0 vn0 avss ibg_200n vn0 vbg_1v2 vp1 avss vbg_1v2 vstart isrc_sel_b vbg_1v2 vstart
+ vp vbg_1v2 avss vn0 vn1 vbg_1v2 vbg_1v2 vp vn0 vstart vbg_1v2 vstart ena vbg_1v2
+ vbg_1v2 sky130_fd_pr__nfet_g5v0d10v5_EC8RE7
Xsky130_fd_pr__pfet_g5v0d10v5_75AJMX_0 avdd avdd avdd vp avdd avdd vp1 avdd avdd vp0
+ vp0 vp1 itest vp avdd vp0 vp0 avdd avdd avdd avdd avdd vp0 avdd vp avdd vp1 vp ibias
+ vn0 sky130_fd_pr__pfet_g5v0d10v5_75AJMX
Xsky130_fd_pr__pfet_g5v0d10v5_Y9J9EP_0 ena avdd avdd isrc_sel_b ena_b isrc_sel avdd
+ avdd sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP
Xsky130_fd_pr__nfet_g5v0d10v5_QZVU2P_1 avss vr ve avss avss vn0 avss vp0 avss ve avss
+ vn0 vn0 vn0 vr vn0 sky130_fd_pr__nfet_g5v0d10v5_QZVU2P
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_4165_119# m1_3409_119# m1_3409_119# m1_5299_7518#
+ m1_1519_7518# m1_385_119# m1_2653_119# m1_385_119# m1_2653_119# m1_6433_119# m1_1897_119#
+ avss m1_6055_7518# m1_3787_7518# m1_2275_7518# m1_1519_7518# m1_6055_7518# m1_4165_119#
+ m1_5299_7518# m1_763_7518# m1_4921_119# m1_763_7518# m1_7189_119# m1_4543_7518#
+ m1_1897_119# m1_7189_119# m1_3031_7518# m1_6811_7518# m1_4921_119# m1_5677_119#
+ m1_5677_119# m1_6811_7518# m1_3031_7518# m1_3787_7518# m1_1141_119# avss m1_4543_7518#
+ m1_1141_119# m1_6433_119# vr m1_2275_7518# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0 vn1 isrc_sel vp avdd vp1 vstart isrc_sel_b
+ ena_b avdd ibg_200n avdd isrc_sel ena_b avdd vp0 vp avdd isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_7JLQGA
Xsky130_fd_pr__nfet_g5v0d10v5_3DCHX4_0 avss avss vn1 avss avss avss avss avss vn1
+ avss avss avss vn1 avss avss avss vn1 vn1 avss vn1 vp1 avss avss avss avss vp1 avss
+ vn1 avss avss avss avss avss vn1 avss vp1 avss vp1 avss vn1 vn1 avss vn1 avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_3DCHX4
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X4 VGND A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_772_151# a_404_1133# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X10 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X11 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X13 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_SCV3UK a_50_n131# a_n50_n157# a_n526_n243# a_n108_n131#
+ a_n266_n131# a_n424_n131# a_208_n131# a_108_n157# a_n208_n157# a_366_n131# a_266_n157#
+ a_n366_n157#
X0 a_n108_n131# a_n208_n157# a_n266_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_208_n131# a_108_n157# a_50_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n266_n131# a_n366_n157# a_n424_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_366_n131# a_266_n157# a_208_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X4 a_50_n131# a_n50_n157# a_n108_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_BZXTE7 a_208_n64# a_n108_n64# a_998_n64# a_n898_n64#
+ a_108_n161# a_50_n64# a_n208_n161# a_266_n161# a_n424_n64# a_524_n64# a_898_n161#
+ a_n366_n161# a_424_n161# a_n998_n161# a_n266_n64# a_366_n64# a_n524_n161# a_582_n161#
+ a_n50_n161# a_840_n64# a_n740_n64# a_n682_n161# a_740_n161# a_682_n64# a_n582_n64#
+ a_n840_n161# w_n1194_n284# a_n1056_n64#
X0 a_n898_n64# a_n998_n161# a_n1056_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_n582_n64# a_n682_n161# a_n740_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_50_n64# a_n50_n161# a_n108_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n740_n64# a_n840_n161# a_n898_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n266_n64# a_n366_n161# a_n424_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n424_n64# a_n524_n161# a_n582_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n108_n64# a_n208_n161# a_n266_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_998_n64# a_898_n161# a_840_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X8 a_682_n64# a_582_n161# a_524_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_840_n64# a_740_n161# a_682_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_366_n64# a_266_n161# a_208_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_524_n64# a_424_n161# a_366_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_208_n64# a_108_n161# a_50_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt schmitt_trigger_ov in out dvdd dvss
Xsky130_fd_pr__nfet_01v8_SCV3UK_1 m out dvss dvss m dvss dvss dvss in out m in sky130_fd_pr__nfet_01v8_SCV3UK
Xsky130_fd_pr__pfet_01v8_BZXTE7_0 dvdd dvdd out m out m in out dvdd dvdd m in dvdd
+ in m m in m out dvdd dvdd in m out m in dvdd dvdd sky130_fd_pr__pfet_01v8_BZXTE7
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GLAJGT m2_n5000_n839# a_3287_n673# a_1629_47#
+ a_1687_21# a_3287_527# a_1687_741# m2_n26_n839# m2_n1684_n839# a_n5003_n673# a_n1629_261#
+ m2_3290_n839# a_n29_n913# a_n1687_n673# a_n3345_n433# a_n1687_47# a_n3287_741# a_1629_n433#
+ a_3345_261# a_n1687_767# a_n29_n193# a_3345_n699# a_3345_n219# a_n3345_287# a_29_261#
+ a_1629_527# a_n5003_527# a_n1629_n939# a_1687_n459# a_n1629_741# a_n3345_n913# a_n29_287#
+ a_1629_n913# a_29_n459# a_n29_47# a_3287_287# a_3345_741# a_29_21# a_n3287_21# m2_4948_n839#
+ a_n29_n673# a_n3345_n193# a_1629_n193# a_n3345_767# a_29_741# a_1687_n939# a_n3287_n459#
+ a_n5003_47# a_1629_287# a_n5003_287# a_n1629_n699# a_n1629_n219# a_n29_767# a_29_n939#
+ a_3287_n433# a_1687_501# a_3287_767# m2_n3342_n839# a_n5003_n433# a_n3345_n673#
+ a_n1629_21# a_n3287_501# a_1629_n673# a_n1687_n433# a_n1687_527# a_n5137_n1073#
+ m2_1632_n839# a_n3287_n939# a_3345_n459# a_1629_767# a_n5003_767# a_1687_n699# a_1687_n219#
+ a_3345_21# a_3287_n913# a_n5003_n913# a_3287_47# a_n3345_47# a_n1629_501# a_n1687_n913#
+ a_29_n699# a_29_n219# a_1687_261# a_3345_501# a_3287_n193# a_n5003_n193# a_n29_n433#
+ a_n3287_261# a_3345_n939# a_n1687_n193# a_n1687_287# a_n3345_527# a_29_501# a_n3287_n699#
+ a_n3287_n219# a_n1629_n459# a_n29_527#
X0 a_n1687_527# a_n3287_501# a_n3345_527# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X1 a_1629_47# a_29_21# a_n29_47# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X2 a_1629_n913# a_29_n939# a_n29_n913# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X3 a_1629_n193# a_29_n219# a_n29_n193# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X4 a_n3345_n433# a_n5003_n433# a_n5003_n433# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X5 a_n1687_287# a_n3287_261# a_n3345_287# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X6 a_3287_n433# a_1687_n459# a_1629_n433# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X7 a_1629_n673# a_29_n699# a_n29_n673# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X8 a_n3345_n913# a_n5003_n913# a_n5003_n913# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X9 a_n1687_767# a_n3287_741# a_n3345_767# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X10 a_n3345_n193# a_n5003_n193# a_n5003_n193# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X11 a_n1687_n433# a_n3287_n459# a_n3345_n433# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X12 a_n29_527# a_n1629_501# a_n1687_527# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X13 a_n1687_47# a_n3287_21# a_n3345_47# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X14 a_3345_21# a_3345_21# a_3287_47# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X15 a_3287_n193# a_1687_n219# a_1629_n193# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X16 a_3287_n913# a_1687_n939# a_1629_n913# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X17 a_n1687_n193# a_n3287_n219# a_n3345_n193# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X18 a_n3345_n673# a_n5003_n673# a_n5003_n673# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X19 a_n1687_n913# a_n3287_n939# a_n3345_n913# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X20 a_n29_287# a_n1629_261# a_n1687_287# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X21 a_3287_n673# a_1687_n699# a_1629_n673# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X22 a_n3345_527# a_n5003_527# a_n5003_527# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X23 a_n1687_n673# a_n3287_n699# a_n3345_n673# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X24 a_n29_767# a_n1629_741# a_n1687_767# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X25 a_3345_n459# a_3345_n459# a_3287_n433# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X26 a_n3345_287# a_n5003_287# a_n5003_287# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X27 a_3345_n219# a_3345_n219# a_3287_n193# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X28 a_3345_n939# a_3345_n939# a_3287_n913# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X29 a_n3345_767# a_n5003_767# a_n5003_767# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X30 a_n3345_47# a_n5003_47# a_n5003_47# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X31 a_1629_527# a_29_501# a_n29_527# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X32 a_3345_n699# a_3345_n699# a_3287_n673# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X33 a_3287_527# a_1687_501# a_1629_527# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X34 a_1629_287# a_29_261# a_n29_287# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X35 a_3345_501# a_3345_501# a_3287_527# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X36 a_3287_287# a_1687_261# a_1629_287# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X37 a_n29_47# a_n1629_21# a_n1687_47# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X38 a_1629_767# a_29_741# a_n29_767# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X39 a_n29_n433# a_n1629_n459# a_n1687_n433# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X40 a_3287_47# a_1687_21# a_1629_47# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X41 a_3287_767# a_1687_741# a_1629_767# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X42 a_3345_261# a_3345_261# a_3287_287# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X43 a_n29_n193# a_n1629_n219# a_n1687_n193# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X44 a_n29_n913# a_n1629_n939# a_n1687_n913# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X45 a_3345_741# a_3345_741# a_3287_767# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X46 a_n29_n673# a_n1629_n699# a_n1687_n673# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X47 a_1629_n433# a_29_n459# a_n29_n433# a_n5137_n1073# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4 a_n100_n344# a_n158_118# a_n100_21# a_100_n612#
+ a_100_483# a_n100_n709# a_100_n247# a_n158_n612# a_n100_386# a_n158_n247# a_100_118#
+ w_n358_n909# a_n158_483#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_483# a_n100_386# a_n158_483# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n247# a_n100_n344# a_n158_n247# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n612# a_n100_n709# a_n158_n612# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3HV7M9 a_3345_n161# a_n1687_n64# a_n1629_n161#
+ a_n4945_n161# w_n5203_n362# a_1687_n161# a_n3345_n64# a_29_n161# a_3287_n64# a_n29_n64#
+ a_n3287_n161# a_1629_n64# a_n5003_n64# a_4945_n64#
X0 a_n29_n64# a_n1629_n161# a_n1687_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n3345_n64# a_n4945_n161# a_n5003_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2 a_1629_n64# a_29_n161# a_n29_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_3287_n64# a_1687_n161# a_1629_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_4945_n64# a_3345_n161# a_3287_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X5 a_n1687_n64# a_n3287_n161# a_n3345_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T82T27 a_1629_47# a_1687_21# a_n1687_47# a_4945_n309#
+ a_n1629_n335# a_n5137_n469# a_n4945_n335# a_n29_47# a_29_21# a_n3287_21# a_1687_n335#
+ a_3287_n309# a_n5003_n309# a_29_n335# a_n1687_n309# a_n5003_47# a_n4945_21# a_n3287_n335#
+ a_n1629_21# a_3345_21# a_n29_n309# a_3287_47# a_n3345_47# a_3345_n335# a_n3345_n309#
+ a_1629_n309# a_4945_47#
X0 a_1629_47# a_29_21# a_n29_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n1687_47# a_n3287_21# a_n3345_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 a_4945_47# a_3345_21# a_3287_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X3 a_1629_n309# a_29_n335# a_n29_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_n3345_n309# a_n4945_n335# a_n5003_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X5 a_3287_n309# a_1687_n335# a_1629_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n1687_n309# a_n3287_n335# a_n3345_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n3345_47# a_n4945_21# a_n5003_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X8 a_n29_47# a_n1629_21# a_n1687_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_4945_n309# a_3345_n335# a_3287_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X10 a_3287_47# a_1687_21# a_1629_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_n29_n309# a_n1629_n335# a_n1687_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z a_n100_199# a_100_n487# a_100_581# a_100_n131#
+ a_n158_n487# a_n100_n157# a_n100_555# a_100_n843# a_n158_n131# a_n158_225# a_n100_n869#
+ a_n158_581# a_n158_n843# a_n100_n513# a_n292_n1003# a_100_225#
X0 a_100_n131# a_n100_n157# a_n158_n131# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_581# a_n100_555# a_n158_581# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n843# a_n100_n869# a_n158_n843# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_225# a_n100_199# a_n158_225# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n487# a_n100_n513# a_n158_n487# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8FRRWQ a_n5003_n7# a_n29_n1003# a_3345_n602#
+ a_3345_n851# a_n3345_740# a_4945_n256# a_1629_n1003# a_n4945_n1100# a_n5003_989#
+ a_n5003_242# a_1629_989# a_1629_242# a_n1629_n104# a_n3345_n505# a_n5003_491# a_1629_491#
+ a_n1629_n353# a_1687_145# a_n3345_n754# a_1687_394# a_1629_n505# a_1629_n754# a_n29_740#
+ a_3287_740# a_4945_242# a_4945_989# a_n3287_145# a_n3287_394# a_4945_491# a_n1629_n1100#
+ a_3287_n1003# a_n4945_n104# a_n3345_n7# a_3287_n7# a_n4945_n353# a_4945_n505# a_4945_n754#
+ a_1687_n104# a_3287_n256# a_1687_n353# a_1629_740# a_n1629_145# a_n5003_n256# a_n1629_n602#
+ a_n5003_740# a_n1629_394# a_n1629_n851# a_1687_643# a_1687_892# a_n1687_n256# a_n5003_n1003#
+ a_3345_145# a_29_n104# w_n5203_n1300# a_4945_740# a_n4945_145# a_n3287_n1100# a_n3287_643#
+ a_3345_394# a_29_n353# a_n4945_394# a_n3287_892# a_3345_n1100# a_n3345_n1003# a_29_145#
+ a_4945_n7# a_29_394# a_n4945_n602# a_n1687_989# a_n1687_242# a_n4945_n851# a_n1687_491#
+ a_n3287_n104# a_1629_n7# a_n3287_n353# a_1687_n1100# a_n1687_n1003# a_1687_n602#
+ a_3287_n505# a_n5003_n505# a_n1687_n7# a_1687_n851# a_3287_n754# a_n5003_n754# a_n1629_643#
+ a_n1629_892# a_n1687_n505# a_n1687_n754# a_n29_n256# a_29_n602# a_3345_643# a_29_n851#
+ a_n4945_643# a_3345_892# a_n4945_892# a_29_643# a_29_892# a_n1687_740# a_29_n1100#
+ a_n3287_n602# a_3345_n104# a_n3287_n851# a_n3345_242# a_3345_n353# a_n3345_989#
+ a_n29_n7# a_n3345_491# a_n3345_n256# a_n29_n505# a_1629_n256# a_n29_n754# a_n29_989#
+ a_n29_242# a_3287_989# a_n29_491# a_3287_242# a_4945_n1003# a_3287_491#
X0 a_n1687_n7# a_n3287_n104# a_n3345_n7# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X1 a_4945_n7# a_3345_n104# a_3287_n7# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X2 a_1629_n256# a_29_n353# a_n29_n256# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X3 a_4945_740# a_3345_643# a_3287_740# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X4 a_n3345_n1003# a_n4945_n1100# a_n5003_n1003# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X5 a_n3345_n256# a_n4945_n353# a_n5003_n256# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X6 a_1629_989# a_29_892# a_n29_989# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X7 a_n1687_491# a_n3287_394# a_n3345_491# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X8 a_1629_242# a_29_145# a_n29_242# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X9 a_3287_n256# a_1687_n353# a_1629_n256# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X10 a_3287_989# a_1687_892# a_1629_989# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X11 a_3287_242# a_1687_145# a_1629_242# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X12 a_n1687_n256# a_n3287_n353# a_n3345_n256# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X13 a_4945_n754# a_3345_n851# a_3287_n754# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X14 a_n1687_n1003# a_n3287_n1100# a_n3345_n1003# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X15 a_4945_n1003# a_3345_n1100# a_3287_n1003# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X16 a_4945_989# a_3345_892# a_3287_989# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X17 a_4945_242# a_3345_145# a_3287_242# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X18 a_1629_n505# a_29_n602# a_n29_n505# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X19 a_1629_n1003# a_29_n1100# a_n29_n1003# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X20 a_n29_491# a_n1629_394# a_n1687_491# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X21 a_n3345_n7# a_n4945_n104# a_n5003_n7# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X22 a_n3345_n505# a_n4945_n602# a_n5003_n505# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X23 a_n1687_740# a_n3287_643# a_n3345_740# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X24 a_4945_n256# a_3345_n353# a_3287_n256# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X25 a_3287_n1003# a_1687_n1100# a_1629_n1003# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X26 a_3287_n505# a_1687_n602# a_1629_n505# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X27 a_n3345_491# a_n4945_394# a_n5003_491# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X28 a_n29_n7# a_n1629_n104# a_n1687_n7# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X29 a_n1687_n505# a_n3287_n602# a_n3345_n505# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X30 a_n29_n754# a_n1629_n851# a_n1687_n754# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X31 a_3287_n7# a_1687_n104# a_1629_n7# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X32 a_n29_740# a_n1629_643# a_n1687_740# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X33 a_n1687_989# a_n3287_892# a_n3345_989# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X34 a_n1687_242# a_n3287_145# a_n3345_242# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X35 a_1629_491# a_29_394# a_n29_491# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X36 a_n29_n256# a_n1629_n353# a_n1687_n256# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X37 a_4945_n505# a_3345_n602# a_3287_n505# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X38 a_3287_491# a_1687_394# a_1629_491# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X39 a_n29_n1003# a_n1629_n1100# a_n1687_n1003# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X40 a_n3345_740# a_n4945_643# a_n5003_740# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X41 a_4945_491# a_3345_394# a_3287_491# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=8
X42 a_n29_989# a_n1629_892# a_n1687_989# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X43 a_n29_242# a_n1629_145# a_n1687_242# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X44 a_1629_n754# a_29_n851# a_n29_n754# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X45 a_1629_n7# a_29_n104# a_n29_n7# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X46 a_n3345_n754# a_n4945_n851# a_n5003_n754# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X47 a_1629_740# a_29_643# a_n29_740# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X48 a_3287_n754# a_1687_n851# a_1629_n754# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X49 a_n3345_989# a_n4945_892# a_n5003_989# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X50 a_3287_740# a_1687_643# a_1629_740# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X51 a_n3345_242# a_n4945_145# a_n5003_242# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=8
X52 a_n29_n505# a_n1629_n602# a_n1687_n505# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
X53 a_n1687_n754# a_n3287_n851# a_n3345_n754# w_n5203_n1300# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z a_861_n131# a_207_n157# a_n861_n157# a_n563_n131#
+ a_683_n131# a_n919_n131# a_29_n157# a_n683_n157# a_n385_n131# a_n1053_n291# a_741_n157#
+ a_505_n131# a_n505_n157# a_563_n157# a_n207_n131# a_327_n131# a_n327_n157# a_385_n157#
+ a_n29_n131# a_149_n131# a_n741_n131# a_n149_n157#
X0 a_n563_n131# a_n683_n157# a_n741_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1 a_505_n131# a_385_n157# a_327_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2 a_n385_n131# a_n505_n157# a_n563_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X3 a_327_n131# a_207_n157# a_149_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X4 a_149_n131# a_29_n157# a_n29_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X5 a_861_n131# a_741_n157# a_683_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X6 a_n207_n131# a_n327_n157# a_n385_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X7 a_n741_n131# a_n861_n157# a_n919_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X8 a_683_n131# a_563_n157# a_505_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X9 a_n29_n131# a_n149_n157# a_n207_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_W8MWAU a_n741_n136# w_n1119_n362# a_861_n136#
+ a_n327_n162# a_385_n162# a_n563_n136# a_683_n136# a_n149_n162# a_n919_n136# a_207_n162#
+ a_n385_n136# a_n861_n162# a_505_n136# a_29_n162# a_n207_n136# a_n683_n162# a_741_n162#
+ a_327_n136# a_n505_n162# a_n29_n136# a_563_n162# a_149_n136#
X0 a_861_n136# a_741_n162# a_683_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X1 a_n207_n136# a_n327_n162# a_n385_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2 a_n741_n136# a_n861_n162# a_n919_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 a_683_n136# a_563_n162# a_505_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X4 a_n29_n136# a_n149_n162# a_n207_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X5 a_n563_n136# a_n683_n162# a_n741_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X6 a_505_n136# a_385_n162# a_327_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X7 a_n385_n136# a_n505_n162# a_n563_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X8 a_327_n136# a_207_n162# a_149_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X9 a_149_n136# a_29_n162# a_n29_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
.ends

.subckt comparator_ov ibias out ena vinn vinp vt avdd
Xsky130_fd_pr__nfet_g5v0d10v5_GLAJGT_1 vt vnn vt vinn vnn vinn vpp vt vt vinp vnn
+ vpp vt vnn vt vinn vt vt vt vpp vt vt vnn vinp vt vt vinp vinn vinp vnn vpp vt vinp
+ vpp vnn vt vinp vinn vt vpp vnn vt vnn vinp vinn vinn vt vt vt vinp vinp vpp vinp
+ vnn vinn vnn vnn vt vnn vinp vinn vt vt vt vt vt vinn vt vt vt vinn vinn vt vnn
+ vt vnn vnn vinp vt vinp vinp vinn vt vnn vt vpp vinn vt vt vt vnn vinp vinn vinn
+ vinp vpp sky130_fd_pr__nfet_g5v0d10v5_GLAJGT
Xsky130_fd_pr__pfet_g5v0d10v5_5H9LZ4_0 ena avdd ena vn vpp ena_b ena_b ibias ena avdd
+ vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4
Xsky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0 avdd vm vnn avdd avdd vpp avdd vpp avdd avdd
+ vnn n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5_3HV7M9
Xsky130_fd_pr__nfet_g5v0d10v5_T82T27_1 n0 vm vm vt vn vt vt vt vm vm vn vt vt vn vn
+ vt vt vn vm vt vt vt vt vt vt vt vt sky130_fd_pr__nfet_g5v0d10v5_T82T27
Xsky130_fd_pr__nfet_g5v0d10v5_GG9S2Z_0 ena vm vn vn vt ena_b ena n0 vt vt ena_b ibias
+ vt ena_b vt ena_b sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z
Xsky130_fd_pr__pfet_g5v0d10v5_8FRRWQ_0 avdd avdd avdd avdd avdd avdd vnn avdd avdd
+ avdd vnn vnn vnn avdd avdd vnn vnn vnn avdd vnn vnn vnn avdd avdd avdd avdd vpp
+ vpp avdd vnn avdd avdd avdd avdd avdd avdd avdd vpp avdd vpp vnn vpp avdd vnn avdd
+ vpp vnn vnn vnn vpp avdd avdd vpp avdd avdd avdd vnn vpp avdd vpp avdd vpp avdd
+ avdd vnn avdd vnn avdd vpp vpp avdd vpp vnn vnn vnn vpp vpp vpp avdd avdd vpp vpp
+ avdd avdd vpp vpp vpp vpp avdd vpp avdd vpp avdd avdd avdd vnn vnn vpp vpp vnn avdd
+ vnn avdd avdd avdd avdd avdd avdd avdd vnn avdd avdd avdd avdd avdd avdd avdd avdd
+ sky130_fd_pr__pfet_g5v0d10v5_8FRRWQ
Xsky130_fd_pr__nfet_g5v0d10v5_HZHY2Z_0 vt n1 n1 vt n1 vt n1 n1 out vt n0 vt n1 n0
+ vt out n1 n1 out vt out n1 sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z
Xsky130_fd_pr__pfet_g5v0d10v5_W8MWAU_0 out avdd avdd n1 n1 avdd n1 n1 avdd n1 out
+ n1 avdd n1 avdd n1 n0 out n1 out n0 avdd sky130_fd_pr__pfet_g5v0d10v5_W8MWAU
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LUWKLG c2_n3269_n19000# m4_n3349_n19080#
X0 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X3 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X4 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X5 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 Base Collector Emitter m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544
.ends

.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt overvoltage_ana otrip_decoded[14] otrip_decoded[13] otrip_decoded[11] otrip_decoded[10]
+ otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[3] otrip_decoded[1]
+ otrip_decoded[0] ena dvdd isrc_sel itest ibg_200n ovout vin otrip_decoded[4] vbg_1v2
+ otrip_decoded[8] otrip_decoded[2] avdd otrip_decoded[15] otrip_decoded[9] otrip_decoded[12]
+ avss ibias_gen_ov_0/ve dvss
Xsky130_fd_sc_hvl__lsbufhv2lv_1_0 dcomp dvdd dvss dvss avdd avdd vl sky130_fd_sc_hvl__lsbufhv2lv_1
Xrstring_mux_ov_0 vin ibias_gen_ov_0/ena sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/X sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/X
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/X sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/X
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/X sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/X
+ rstring_mux_ov_0/otrip_decoded_avdd[9] rstring_mux_ov_0/otrip_decoded_avdd[8] rstring_mux_ov_0/otrip_decoded_avdd[7]
+ rstring_mux_ov_0/otrip_decoded_avdd[6] rstring_mux_ov_0/otrip_decoded_avdd[5] rstring_mux_ov_0/otrip_decoded_avdd[4]
+ rstring_mux_ov_0/otrip_decoded_avdd[3] rstring_mux_ov_0/otrip_decoded_avdd[2] rstring_mux_ov_0/otrip_decoded_avdd[1]
+ rstring_mux_ov_0/otrip_decoded_avdd[0] rstring_mux_ov_0/vtop avdd avss rstring_mux_ov
Xibias_gen_ov_0 itest ibias_gen_ov_0/ibias ibg_200n vbg_1v2 ibias_gen_ov_0/isrc_sel
+ ibias_gen_ov_0/ena ibias_gen_ov_0/ve avss avdd ibias_gen_ov
Xsky130_fd_sc_hd__inv_4_0 schmitt_trigger_ov_0/out dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_0/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] otrip_decoded[0] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] otrip_decoded[1] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] otrip_decoded[2] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] otrip_decoded[3] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2] otrip_decoded[4] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2] otrip_decoded[5] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3] otrip_decoded[6] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3] otrip_decoded[7] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4] otrip_decoded[8] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[8]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4] otrip_decoded[9] dvdd dvss dvss avdd avdd rstring_mux_ov_0/otrip_decoded_avdd[9]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5] otrip_decoded[10] dvdd dvss dvss avdd avdd
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5]/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5] otrip_decoded[11] dvdd dvss dvss avdd avdd
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5]/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6] otrip_decoded[12] dvdd dvss dvss avdd avdd
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6]/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6] otrip_decoded[13] dvdd dvss dvss avdd avdd
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6]/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7] otrip_decoded[14] dvdd dvss dvss avdd avdd
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7]/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7] otrip_decoded[15] dvdd dvss dvss avdd avdd
+ sky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7]/X sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8] ena dvdd dvss dvss avdd avdd ibias_gen_ov_0/ena
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8] isrc_sel dvdd dvss dvss avdd avdd ibias_gen_ov_0/isrc_sel
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xschmitt_trigger_ov_0 schmitt_trigger_ov_0/in schmitt_trigger_ov_0/out dvdd dvss schmitt_trigger_ov
Xcomparator_ov_0 ibias_gen_ov_0/ibias dcomp ibias_gen_ov_0/ena vbg_1v2 vin avss avdd
+ comparator_ov
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_n11325_2001# m1_n11325_2001# m1_n12081_2001#
+ m1_n10191_9400# m1_n13971_9400# m1_n14349_2001# m1_n12081_2001# vl m1_n12837_2001#
+ m1_n8301_2001# m1_n12837_2001# avss m1_n9435_9400# m1_n10947_9400# m1_n13215_9400#
+ m1_n13215_9400# m1_n8679_9400# m1_n10569_2001# m1_n9435_9400# m1_n13971_9400# m1_n10569_2001#
+ m1_n14727_9400# m1_n8301_2001# m1_n10947_9400# m1_n13593_2001# schmitt_trigger_ov_0/in
+ m1_n11703_9400# m1_n8679_9400# m1_n9813_2001# m1_n9057_2001# m1_n9813_2001# m1_n7923_9400#
+ m1_n12459_9400# m1_n11703_9400# m1_n13593_2001# m1_n14727_9400# m1_n10191_9400#
+ m1_n14349_2001# m1_n9057_2001# m1_n7923_9400# m1_n12459_9400# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 schmitt_trigger_ov_0/in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xsky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 avss avss ibias_gen_ov_0/ve sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 m=1
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_4_0/Y dvss dvss dvdd dvdd ovout sky130_fd_sc_hd__inv_16
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
X0 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_91_199# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6 a_245_297# C a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_341_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X8 a_91_199# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X9 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt overvoltage_dig otrip_decoded[15] otrip_decoded[14] otrip_decoded[13] otrip_decoded[12]
+ otrip_decoded[11] otrip_decoded[10] otrip_decoded[9] otrip_decoded[8] otrip_decoded[7]
+ otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3] otrip_decoded[2]
+ otrip_decoded[1] otrip_decoded[0] otrip[3] otrip[2] otrip[1] otrip[0] VPWR VGND
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput20 net20 VGND VGND VPWR VPWR otrip_decoded[9] sky130_fd_sc_hd__buf_2
Xoutput7 net7 VGND VGND VPWR VPWR otrip_decoded[11] sky130_fd_sc_hd__buf_2
XFILLER_0_13_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput10 net10 VGND VGND VPWR VPWR otrip_decoded[14] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR otrip_decoded[12] sky130_fd_sc_hd__buf_2
XFILLER_0_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR otrip_decoded[13] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR otrip_decoded[15] sky130_fd_sc_hd__buf_2
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_4_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
X_09_ net25 net23 net22 net28 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08_ net28 net26 net24 net22 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__nor4b_1
XFILLER_0_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07_ net21 net27 net26 net24 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and4b_1
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06_ net21 net27 net25 net23 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and4bb_1
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[8] sky130_fd_sc_hd__buf_2
X_05_ net21 net25 net23 net27 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and4bb_1
XFILLER_0_13_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout21 net4 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_04_ net21 net27 net25 net23 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor4b_1
XFILLER_0_2_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout22 net4 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 otrip[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_03_ net21 net23 net25 net27 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout23 net3 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 otrip[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_02_ net21 net27 net23 net25 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor4b_1
XFILLER_0_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout24 net3 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
X_01_ net21 net25 net23 net27 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor4b_1
Xinput3 otrip[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout25 net2 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 otrip[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_00_ net21 net27 net25 net23 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__nor4_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout26 net2 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout27 net1 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout28 net1 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ net22 net28 net26 net24 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__and4_1
XFILLER_0_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14_ net28 net26 net24 net22 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__and4b_1
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13_ net26 net24 net22 net28 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12_ net27 net25 net23 net21 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11_ net24 net26 net28 net22 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__and4b_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10_ net27 net23 net25 net21 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput6 net6 VGND VGND VPWR VPWR otrip_decoded[10] sky130_fd_sc_hd__buf_2
.ends

.subckt sky130_fd_pr__nfet_01v8_D5N54F a_n287_n188# a_761_n100# a_819_n188# a_n29_n100#
+ a_345_n188# a_n919_n188# a_n445_n188# a_n1079_n274# a_n187_n100# a_503_n188# a_n819_n100#
+ a_n603_n188# a_n345_n100# a_661_n188# a_n977_n100# a_n761_n188# a_129_n100# a_n503_n100#
+ a_n661_n100# a_287_n100# a_919_n100# a_445_n100# a_29_n188# a_n129_n188# a_603_n100#
+ a_187_n188#
X0 a_287_n100# a_187_n188# a_129_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_919_n100# a_819_n188# a_761_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X2 a_445_n100# a_345_n188# a_287_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_603_n100# a_503_n188# a_445_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n661_n100# a_n761_n188# a_n819_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_129_n100# a_29_n188# a_n29_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n187_n100# a_n287_n188# a_n345_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n819_n100# a_n919_n188# a_n977_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X8 a_n345_n100# a_n445_n188# a_n503_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n503_n100# a_n603_n188# a_n661_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_n29_n100# a_n129_n188# a_n187_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_761_n100# a_661_n188# a_603_n100# a_n1079_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_53744R a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_ajc_ip__overvoltage avdd dvdd vbg_1v2 ovout itest otrip[3] otrip[2]
+ otrip[1] otrip[0] vin ena isrc_sel ibg_200n avss dvss
Xovervoltage_ana_0 overvoltage_dig_0/otrip_decoded[14] overvoltage_dig_0/otrip_decoded[13]
+ overvoltage_dig_0/otrip_decoded[11] overvoltage_dig_0/otrip_decoded[10] overvoltage_dig_0/otrip_decoded[7]
+ overvoltage_dig_0/otrip_decoded[6] overvoltage_dig_0/otrip_decoded[5] overvoltage_dig_0/otrip_decoded[3]
+ overvoltage_dig_0/otrip_decoded[1] overvoltage_dig_0/otrip_decoded[0] ena dvdd isrc_sel
+ itest ibg_200n ovout vin overvoltage_dig_0/otrip_decoded[4] vbg_1v2 overvoltage_dig_0/otrip_decoded[8]
+ overvoltage_dig_0/otrip_decoded[2] avdd overvoltage_dig_0/otrip_decoded[15] overvoltage_dig_0/otrip_decoded[9]
+ overvoltage_dig_0/otrip_decoded[12] avss overvoltage_ana_0/ibias_gen_ov_0/ve dvss
+ overvoltage_ana
Xovervoltage_dig_0 overvoltage_dig_0/otrip_decoded[15] overvoltage_dig_0/otrip_decoded[14]
+ overvoltage_dig_0/otrip_decoded[13] overvoltage_dig_0/otrip_decoded[12] overvoltage_dig_0/otrip_decoded[11]
+ overvoltage_dig_0/otrip_decoded[10] overvoltage_dig_0/otrip_decoded[9] overvoltage_dig_0/otrip_decoded[8]
+ overvoltage_dig_0/otrip_decoded[7] overvoltage_dig_0/otrip_decoded[6] overvoltage_dig_0/otrip_decoded[5]
+ overvoltage_dig_0/otrip_decoded[4] overvoltage_dig_0/otrip_decoded[3] overvoltage_dig_0/otrip_decoded[2]
+ overvoltage_dig_0/otrip_decoded[1] overvoltage_dig_0/otrip_decoded[0] otrip[3] otrip[2]
+ otrip[1] otrip[0] dvdd dvss overvoltage_dig
Xsky130_fd_pr__nfet_01v8_D5N54F_0 dvss ena dvss dvss dvss dvss dvss dvss otrip[1]
+ dvss otrip[3] dvss dvss dvss dvss dvss otrip[0] otrip[2] dvss dvss dvss isrc_sel
+ dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_D5N54F
Xsky130_fd_pr__nfet_01v8_53744R_0 dvss vin dvss dvss sky130_fd_pr__nfet_01v8_53744R
Xsky130_fd_pr__nfet_01v8_53744R_1 dvss vbg_1v2 dvss dvss sky130_fd_pr__nfet_01v8_53744R
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PXF6AN a_1235_n100# a_n287_n188# a_761_n100#
+ a_819_n188# a_n1077_n188# a_n29_n100# a_345_n188# a_n919_n188# a_977_n188# a_n445_n188#
+ a_n187_n100# a_n1235_n188# a_503_n188# a_n819_n100# a_n603_n188# a_n345_n100# a_1135_n188#
+ a_661_n188# a_n977_n100# a_n1135_n100# a_n761_n188# a_129_n100# a_n503_n100# a_n1293_n100#
+ a_n661_n100# a_287_n100# a_919_n100# a_445_n100# a_1077_n100# a_29_n188# a_n1427_n322#
+ a_n129_n188# a_603_n100# a_187_n188#
X0 a_919_n100# a_819_n188# a_761_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_445_n100# a_345_n188# a_287_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_603_n100# a_503_n188# a_445_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n977_n100# a_n1077_n188# a_n1135_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n1135_n100# a_n1235_n188# a_n1293_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X5 a_n661_n100# a_n761_n188# a_n819_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_129_n100# a_29_n188# a_n29_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n187_n100# a_n287_n188# a_n345_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_n819_n100# a_n919_n188# a_n977_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n345_n100# a_n445_n188# a_n503_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_n503_n100# a_n603_n188# a_n661_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_n29_n100# a_n129_n188# a_n187_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_1077_n100# a_977_n188# a_919_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_761_n100# a_661_n188# a_603_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_287_n100# a_187_n188# a_129_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_1235_n100# a_1135_n188# a_1077_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt brownout_dig VPWR brout_filt dcomp ena force_dis_rc_osc force_ena_rc_osc force_short_oneshot
+ osc_ck otrip[0] otrip[1] otrip[2] vtrip[0] vtrip[1] vtrip[2] osc_ena otrip_decoded[0]
+ otrip_decoded[1] otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6]
+ otrip_decoded[7] outb_unbuf timed_out vtrip_decoded[0] vtrip_decoded[1] vtrip_decoded[2]
+ vtrip_decoded[3] vtrip_decoded[4] vtrip_decoded[5] vtrip_decoded[6] vtrip_decoded[7]
+ otrip_decoded[2] VGND
XFILLER_0_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_062_ net9 net7 net8 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and3_1
X_114_ clknet_1_1__leaf_osc_ck _010_ net3 VGND VGND VPWR VPWR cnt\[8\] sky130_fd_sc_hd__dfstp_1
X_045_ net1 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
Xoutput31 net31 VGND VGND VPWR VPWR vtrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_061_ net7 net8 net9 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and3b_1
X_044_ net4 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
X_113_ clknet_1_1__leaf_osc_ck _009_ net33 VGND VGND VPWR VPWR cnt\[7\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_13_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ net8 net7 net9 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and3b_1
X_043_ net32 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_112_ clknet_1_0__leaf_osc_ck _008_ net33 VGND VGND VPWR VPWR cnt\[6\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR outb_unbuf sky130_fd_sc_hd__buf_2
XFILLER_0_13_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_111_ clknet_1_0__leaf_osc_ck _007_ net33 VGND VGND VPWR VPWR cnt\[5\] sky130_fd_sc_hd__dfstp_1
Xoutput23 net23 VGND VGND VPWR VPWR timed_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ clknet_1_0__leaf_osc_ck _006_ net33 VGND VGND VPWR VPWR cnt\[4\] sky130_fd_sc_hd__dfstp_1
Xoutput24 net24 VGND VGND VPWR VPWR vtrip_decoded[0] sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
XFILLER_0_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput25 net25 VGND VGND VPWR VPWR vtrip_decoded[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
X_099_ cnt\[9\] _022_ cnt\[10\] VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a21o_1
Xoutput26 net26 VGND VGND VPWR VPWR vtrip_decoded[2] sky130_fd_sc_hd__clkbuf_4
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_119__35 VGND VGND VPWR VPWR net35 _119__35/LO sky130_fd_sc_hd__conb_1
X_098_ net23 _023_ _028_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_7_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput27 net27 VGND VGND VPWR VPWR vtrip_decoded[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
X_097_ cnt\[9\] _022_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__xor2_1
Xoutput28 net28 VGND VGND VPWR VPWR vtrip_decoded[4] sky130_fd_sc_hd__clkbuf_4
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_096_ cnt\[8\] _035_ net6 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR vtrip_decoded[5] sky130_fd_sc_hd__clkbuf_4
X_079_ cnt\[2\] _030_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
X_095_ _038_ _021_ net38 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_078_ _038_ _040_ net32 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a21oi_1
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout32 clr_cnt VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
X_094_ cnt\[8\] _035_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__xnor2_1
X_077_ _030_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout33 net3 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
X_093_ _038_ _020_ net32 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21oi_1
X_076_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 brout_filt VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ net7 net8 net9 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__nor3b_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 dcomp VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_092_ cnt\[7\] _034_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__xor2_1
X_075_ net39 _038_ net32 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a21oi_1
X_058_ net9 net7 net8 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3b_1
XFILLER_0_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput3 ena VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_074_ net6 net23 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nor2_2
X_091_ _038_ _019_ net32 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21oi_1
X_057_ net9 net7 net8 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_109_ clknet_1_0__leaf_osc_ck _005_ net33 VGND VGND VPWR VPWR cnt\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ _034_ _018_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand2_1
Xinput4 force_dis_rc_osc VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_073_ net2 net33 VGND VGND VPWR VPWR dcomp_ena_rsb sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_6_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_056_ net9 net8 net7 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
X_108_ clknet_1_1__leaf_osc_ck _004_ net33 VGND VGND VPWR VPWR cnt\[2\] sky130_fd_sc_hd__dfstp_1
Xinput5 force_ena_rc_osc VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_072_ net33 _029_ _037_ net5 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__a31o_1
X_055_ net9 net7 net8 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__nor3_1
X_107_ clknet_1_0__leaf_osc_ck _003_ net33 VGND VGND VPWR VPWR cnt\[1\] sky130_fd_sc_hd__dfstp_1
X_118__34 VGND VGND VPWR VPWR _118__34/HI net34 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 force_short_oneshot VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_071_ dcomp_retimed net2 net23 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__or3b_1
X_106_ clknet_1_0__leaf_osc_ck _002_ net33 VGND VGND VPWR VPWR cnt\[0\] sky130_fd_sc_hd__dfstp_1
X_054_ dcomp_retimed net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_070_ net12 net11 net10 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__and3_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 otrip[0] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 vtrip[0] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
X_053_ cnt\[8\] cnt\[11\] _035_ _036_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__and4_2
XFILLER_0_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ net1 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
Xinput8 otrip[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 vtrip[1] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
X_104_ net23 _026_ _027_ _028_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_10_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_052_ cnt\[9\] cnt\[10\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and2_1
X_121_ clknet_1_1__leaf_osc_ck net2 dcomp_ena_rsb VGND VGND VPWR VPWR dcomp_retimed
+ sky130_fd_sc_hd__dfrtp_1
Xinput9 otrip[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 vtrip[2] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_051_ cnt\[4\] cnt\[7\] _031_ _033_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and4_1
X_120_ clknet_1_0__leaf_osc_ck net37 _001_ VGND VGND VPWR VPWR clr_cnt_sb sky130_fd_sc_hd__dfrtp_1
X_103_ _036_ _022_ cnt\[11\] VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 clr_cnt_sb VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
X_102_ cnt\[11\] _036_ _022_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and3b_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
X_050_ _032_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand2_1
Xhold2 clr_cnt_sb_stg1 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_101_ _028_ net23 _024_ _025_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 clr_cnt VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _036_ _022_ net32 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a21oi_1
Xhold4 cnt\[0\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_5_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ cnt\[5\] cnt\[4\] _031_ cnt\[6\] VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ _038_ _017_ net32 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_9_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ cnt\[5\] _032_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_086_ _038_ _016_ net32 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a21oi_1
X_069_ net10 net11 net12 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _032_ _015_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__or2_1
X_068_ net11 net10 net12 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__and3b_1
X_067_ net11 net10 net12 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_13_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_084_ cnt\[4\] _031_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nor2_1
X_119_ clknet_1_0__leaf_osc_ck net35 _000_ VGND VGND VPWR VPWR clr_cnt_sb_stg1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_083_ _038_ _014_ net32 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_066_ net12 net11 net10 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__and3b_1
X_118_ clknet_1_0__leaf_osc_ck net34 net36 VGND VGND VPWR VPWR clr_cnt sky130_fd_sc_hd__dfstp_1
X_049_ cnt\[5\] cnt\[6\] VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_4_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_065_ net12 net10 net11 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__nor3b_1
X_082_ _031_ _042_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_117_ clknet_1_1__leaf_osc_ck _013_ net3 VGND VGND VPWR VPWR cnt\[11\] sky130_fd_sc_hd__dfstp_1
X_048_ cnt\[4\] _031_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__and2_1
X_081_ cnt\[1\] cnt\[0\] cnt\[2\] cnt\[3\] VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_064_ net12 net11 net10 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__nor3b_1
X_047_ cnt\[1\] cnt\[0\] cnt\[3\] cnt\[2\] VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and4_1
X_116_ clknet_1_1__leaf_osc_ck _012_ net3 VGND VGND VPWR VPWR cnt\[10\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_063_ net12 net11 net10 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nor3_1
X_080_ _038_ _041_ net32 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_115_ clknet_1_1__leaf_osc_ck _011_ net3 VGND VGND VPWR VPWR cnt\[9\] sky130_fd_sc_hd__dfstp_1
X_046_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput30 net30 VGND VGND VPWR VPWR vtrip_decoded[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_V6EN4F a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XTZQRT a_n287_n188# a_761_n100# a_n29_n100# a_345_n188#
+ a_n953_n322# a_n445_n188# a_n187_n100# a_503_n188# a_n819_n100# a_n603_n188# a_n345_n100#
+ a_661_n188# a_n761_n188# a_129_n100# a_n503_n100# a_n661_n100# a_287_n100# a_445_n100#
+ a_29_n188# a_n129_n188# a_603_n100# a_187_n188#
X0 a_445_n100# a_345_n188# a_287_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_603_n100# a_503_n188# a_445_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n661_n100# a_n761_n188# a_n819_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_129_n100# a_29_n188# a_n29_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n187_n100# a_n287_n188# a_n345_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n345_n100# a_n445_n188# a_n503_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n503_n100# a_n603_n188# a_n661_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n29_n100# a_n129_n188# a_n187_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_761_n100# a_661_n188# a_603_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X9 a_287_n100# a_187_n188# a_129_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2 a_n7134_n3916# a_n8646_3484# a_7230_3484#
+ a_n5244_3484# a_8364_n3916# a_12144_3484# a_n7512_n3916# a_6096_n3916# a_n9024_3484#
+ a_n5244_n3916# a_n12048_n3916# a_8742_n3916# a_6474_n3916# a_n330_n3916# a_n708_n3916#
+ a_n12426_n3916# a_48_n3916# a_n5622_n3916# a_n7890_3484# a_7986_3484# a_n12804_3484#
+ a_4584_3484# a_n2598_3484# a_n3354_n3916# a_n10158_n3916# a_n13182_3484# a_1182_3484#
+ a_6852_n3916# a_n12804_n3916# a_11388_n3916# a_4584_n3916# a_n1086_n3916# a_8364_3484#
+ a_n10536_n3916# a_n3732_n3916# a_n6378_3484# a_11766_n3916# a_4962_n3916# a_n1464_n3916#
+ a_n10914_n3916# a_2694_n3916# a_n1842_n3916# a_n9780_n3916# a_n1842_3484# a_1938_3484#
+ a_48_3484# a_n10536_3484# a_n5622_3484# a_5718_3484# a_9498_3484# a_n2220_3484#
+ a_n7890_n3916# a_2316_3484# a_6096_3484# a_12522_3484# a_9120_n3916# a_n9402_3484#
+ a_n6000_3484# a_n6000_n3916# a_7230_n3916# a_7608_n3916# a_426_n3916# a_4962_3484#
+ a_1560_3484# a_n2976_3484# a_804_n3916# a_n4110_n3916# a_8742_3484# a_n6756_3484#
+ a_5340_3484# a_12144_n3916# a_n3354_3484# a_5340_n3916# a_5718_n3916# a_n13312_n4046#
+ a_n12048_3484# a_10254_3484# a_3072_n3916# a_9120_3484# a_12522_n3916# a_n2220_n3916#
+ a_n7134_3484# a_426_3484# a_10254_n3916# a_3450_n3916# a_3828_n3916# a_12900_n3916#
+ a_n708_3484# a_1182_n3916# a_n8268_n3916# a_10632_n3916# a_n10914_3484# a_2694_3484#
+ a_n11292_3484# a_9498_n3916# a_n8646_n3916# a_n9780_3484# a_1560_n3916# a_1938_n3916#
+ a_9876_3484# a_6474_3484# a_12900_3484# a_n4488_3484# a_3072_3484# a_9876_n3916#
+ a_n1086_3484# a_n6378_n3916# a_11388_3484# a_n8268_3484# a_n13182_n3916# a_n6756_n3916#
+ a_n330_3484# a_7986_n3916# a_n4488_n3916# a_n11292_n3916# a_n4866_n3916# a_n2598_n3916#
+ a_n3732_3484# a_3828_3484# a_n11670_n3916# a_n12426_3484# a_10632_3484# a_n2976_n3916#
+ a_n7512_3484# a_7608_3484# a_804_3484# a_n4110_3484# a_4206_3484# a_4206_n3916#
+ a_11010_3484# a_11010_n3916# a_n11670_3484# a_2316_n3916# a_n9024_n3916# a_6852_3484#
+ a_3450_3484# a_n4866_3484# a_n9402_n3916# a_n1464_3484# a_n10158_3484# a_11766_3484#
X0 a_n9024_3484# a_n9024_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 a_9876_3484# a_9876_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 a_n11670_3484# a_n11670_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X3 a_n330_3484# a_n330_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 a_3072_3484# a_3072_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 a_5718_3484# a_5718_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X6 a_6474_3484# a_6474_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X7 a_8742_3484# a_8742_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X8 a_n11292_3484# a_n11292_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X9 a_n10536_3484# a_n10536_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X10 a_n7890_3484# a_n7890_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X11 a_2316_3484# a_2316_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X12 a_5340_3484# a_5340_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X13 a_n12804_3484# a_n12804_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 a_n6756_3484# a_n6756_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 a_n4488_3484# a_n4488_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X16 a_n1086_3484# a_n1086_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X17 a_12144_3484# a_12144_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X18 a_n5622_3484# a_n5622_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X19 a_n3354_3484# a_n3354_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X20 a_11010_3484# a_11010_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X21 a_6096_3484# a_6096_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X22 a_9498_3484# a_9498_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X23 a_7608_3484# a_7608_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X24 a_8364_3484# a_8364_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X25 a_n13182_3484# a_n13182_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X26 a_n10158_3484# a_n10158_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X27 a_n9780_3484# a_n9780_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X28 a_4206_3484# a_4206_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X29 a_7230_3484# a_7230_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X30 a_n12426_3484# a_n12426_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X31 a_n8646_3484# a_n8646_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X32 a_n6378_3484# a_n6378_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X33 a_n7512_3484# a_n7512_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X34 a_n5244_3484# a_n5244_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X35 a_n2220_3484# a_n2220_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X36 a_1938_3484# a_1938_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X37 a_2694_3484# a_2694_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X38 a_4962_3484# a_4962_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X39 a_1560_3484# a_1560_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X40 a_11766_3484# a_11766_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X41 a_n2976_3484# a_n2976_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X42 a_48_3484# a_48_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X43 a_10632_3484# a_10632_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X44 a_12900_3484# a_12900_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X45 a_n1842_3484# a_n1842_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X46 a_804_3484# a_804_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X47 a_9120_3484# a_9120_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X48 a_n12048_3484# a_n12048_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X49 a_n8268_3484# a_n8268_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X50 a_n7134_3484# a_n7134_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X51 a_n4110_3484# a_n4110_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X52 a_7986_3484# a_7986_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X53 a_n9402_3484# a_n9402_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X54 a_4584_3484# a_4584_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X55 a_n6000_3484# a_n6000_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X56 a_n708_3484# a_n708_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X57 a_1182_3484# a_1182_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X58 a_3828_3484# a_3828_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X59 a_6852_3484# a_6852_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X60 a_11388_3484# a_11388_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X61 a_n2598_3484# a_n2598_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X62 a_3450_3484# a_3450_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X63 a_10254_3484# a_10254_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X64 a_n10914_3484# a_n10914_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X65 a_n4866_3484# a_n4866_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X66 a_12522_3484# a_12522_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X67 a_n3732_3484# a_n3732_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X68 a_n1464_3484# a_n1464_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X69 a_426_3484# a_426_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
.ends

.subckt rstring_mux vout_brout ena otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5]
+ otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1]
+ vtrip_decoded_avdd[7] vtrip_decoded_avdd[6] vtrip_decoded_avdd[5] vtrip_decoded_avdd[4]
+ vtrip_decoded_avdd[3] vtrip_decoded_avdd[2] vtrip_decoded_avdd[1] vtrip_decoded_avdd[0]
+ vout_vunder vtop otrip_decoded_avdd[0] avdd avss
Xsky130_fd_pr__nfet_g5v0d10v5_K8JYEQ_0 vout_brout vtrip_decoded_avdd[0] vout_vunder
+ otrip_decoded_avdd[3] vtrip7 vtrip5 otrip_decoded_avdd[5] otrip_decoded_avdd[1]
+ vout_brout vout_brout avss avss otrip_decoded_avdd[6] vout_brout vout_brout vtrip6
+ vtrip4 vtrip2 vout_brout vtrip_decoded_avdd[3] avss vtrip_decoded_avdd[5] vtrip1
+ vtrip_decoded_avdd[0] vout_vunder vout_brout avss avss avss vtrip_decoded_avdd[2]
+ vtrip_decoded_avdd[6] vtrip_decoded_avdd[4] otrip_decoded_avdd[6] vout_vunder vout_brout
+ vtrip0 vout_vunder vout_vunder vtrip_decoded_avdd[1] vtrip_decoded_avdd[7] vtrip_decoded_avdd[5]
+ otrip_decoded_avdd[4] vout_vunder vout_brout vout_brout otrip_decoded_avdd[2] vtrip_decoded_avdd[4]
+ vtrip_decoded_avdd[2] avss otrip_decoded_avdd[4] otrip_decoded_avdd[0] vtrip3 vtrip_decoded_avdd[6]
+ vout_vunder vtrip7 vtrip4 vtrip2 vout_vunder vout_vunder vout_vunder vtrip_decoded_avdd[1]
+ avss avss avss vtrip5 avss vout_vunder vtrip3 vout_vunder vtrip1 avss avss avss
+ vout_vunder otrip_decoded_avdd[7] vout_brout vout_brout avss vout_brout otrip_decoded_avdd[5]
+ otrip_decoded_avdd[3] otrip_decoded_avdd[1] vtrip0 vout_brout vout_brout vtrip_decoded_avdd[3]
+ vout_brout avss vout_vunder vout_vunder vtrip6 vtrip_decoded_avdd[7] otrip_decoded_avdd[0]
+ vout_vunder otrip_decoded_avdd[7] otrip_decoded_avdd[2] sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ
Xsky130_fd_pr__pfet_g5v0d10v5_4Z8MHY_0 vtrip_decoded_b_avdd[1] vout_brout vtrip0 avdd
+ avdd vout_brout avdd vout_brout avdd vout_vunder vout_vunder vtrip6 vout_vunder
+ avdd avdd avdd avdd vout_brout otrip_decoded_b_avdd[7] vout_vunder avdd vtrip7 vtrip5
+ otrip_decoded_b_avdd[5] vout_brout otrip_decoded_b_avdd[3] vout_brout vout_brout
+ otrip_decoded_b_avdd[1] vout_brout vtrip_decoded_b_avdd[3] vtrip4 vout_brout vtrip2
+ vtrip6 otrip_decoded_b_avdd[0] vtrip_decoded_b_avdd[7] otrip_decoded_b_avdd[7] vtrip1
+ otrip_decoded_b_avdd[2] vtrip_decoded_b_avdd[0] vout_vunder vout_brout otrip_decoded_b_avdd[3]
+ otrip_decoded_b_avdd[1] otrip_decoded_b_avdd[5] vtrip0 avdd vout_vunder vout_brout
+ avdd otrip_decoded_b_avdd[6] vout_vunder vout_vunder avdd vout_vunder vtrip_decoded_b_avdd[3]
+ vtrip_decoded_b_avdd[5] vout_brout vout_brout vtrip_decoded_b_avdd[0] avdd vtrip3
+ avdd avdd vtrip_decoded_b_avdd[2] vtrip4 vtrip7 vtrip_decoded_b_avdd[4] vtrip2 otrip_decoded_b_avdd[6]
+ vout_vunder vtrip_decoded_b_avdd[6] vout_vunder vout_vunder vout_vunder vtrip_decoded_b_avdd[1]
+ vtrip_decoded_b_avdd[5] vtrip5 vout_vunder otrip_decoded_b_avdd[4] vtrip_decoded_b_avdd[7]
+ vtrip3 vtrip1 vout_vunder otrip_decoded_b_avdd[2] vout_vunder otrip_decoded_b_avdd[0]
+ otrip_decoded_b_avdd[4] vtrip_decoded_b_avdd[2] vtrip_decoded_b_avdd[4] vout_brout
+ avdd vtrip_decoded_b_avdd[6] vout_brout vout_brout sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY
Xsky130_fd_pr__pfet_g5v0d10v5_WY4TLZ_0 vtop ena_b ena_b avdd avdd avdd ena_b avdd
+ vtop ena_b ena_b ena_b ena_b vtop ena_b avdd vtop ena_b ena_b avdd avdd ena_b vtop
+ avdd avdd ena_b vtop ena_b ena_b ena_b vtop vtop avdd ena_b sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ
Xsky130_fd_sc_hvl__inv_1_0[0] otrip_decoded_avdd[0] avss avss avdd avdd otrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[1] otrip_decoded_avdd[1] avss avss avdd avdd otrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[2] otrip_decoded_avdd[2] avss avss avdd avdd otrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[3] otrip_decoded_avdd[3] avss avss avdd avdd otrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[4] otrip_decoded_avdd[4] avss avss avdd avdd otrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[5] otrip_decoded_avdd[5] avss avss avdd avdd otrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[6] otrip_decoded_avdd[6] avss avss avdd avdd otrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[7] otrip_decoded_avdd[7] avss avss avdd avdd otrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[8] vtrip_decoded_avdd[0] avss avss avdd avdd vtrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[9] vtrip_decoded_avdd[1] avss avss avdd avdd vtrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[10] vtrip_decoded_avdd[2] avss avss avdd avdd vtrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[11] vtrip_decoded_avdd[3] avss avss avdd avdd vtrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[12] vtrip_decoded_avdd[4] avss avss avdd avdd vtrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[13] vtrip_decoded_avdd[5] avss avss avdd avdd vtrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[14] vtrip_decoded_avdd[6] avss avss avdd avdd vtrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[15] vtrip_decoded_avdd[7] avss avss avdd avdd vtrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_1 ena avss avss avdd avdd ena_b sky130_fd_sc_hvl__inv_1
Xsky130_fd_pr__res_xhigh_po_1p41_9VZRJ2_0 m1_6950_n3340# m1_5060_4059# m1_20936_4059#
+ m1_8840_4059# m1_22070_n3340# m1_26228_4059# m1_6194_n3340# m1_19802_n3340# m1_5060_4059#
+ m1_8462_n3340# m1_1658_n3340# m1_22826_n3340# m1_20558_n3340# vtrip0 m1_12998_n3340#
+ m1_1658_n3340# vtrip0 m1_8462_n3340# m1_5816_4059# m1_21692_4059# m1_1280_4059#
+ m1_18668_4059# m1_11108_4059# m1_10730_n3340# m1_3926_n3340# vtop vtrip3 m1_20558_n3340#
+ m1_902_n3340# m1_25094_n3340# m1_18290_n3340# m1_12998_n3340# m1_22448_4059# m1_3170_n3340#
+ m1_9974_n3340# m1_7328_4059# m1_25850_n3340# m1_19046_n3340# m1_12242_n3340# m1_3170_n3340#
+ m1_16778_n3340# m1_12242_n3340# m1_3926_n3340# m1_11864_4059# vtrip5 vtrip1 m1_3548_4059#
+ m1_8084_4059# m1_19424_4059# m1_23204_4059# m1_11864_4059# m1_6194_n3340# vtrip7
+ m1_20180_4059# m1_26228_4059# m1_22826_n3340# m1_4304_4059# m1_8084_4059# m1_7706_n3340#
+ m1_21314_n3340# m1_21314_n3340# vtrip2 m1_18668_4059# vtrip5 m1_11108_4059# vtrip2
+ m1_9974_n3340# m1_22448_4059# m1_7328_4059# m1_19424_4059# m1_25850_n3340# m1_10352_4059#
+ m1_19046_n3340# m1_19802_n3340# avss m1_2036_4059# m1_23960_4059# m1_16778_n3340#
+ m1_23204_4059# m1_26606_n3340# m1_11486_n3340# m1_6572_4059# vtrip1 m1_24338_n3340#
+ m1_17534_n3340# m1_17534_n3340# m1_26606_n3340# m1_13376_4059# vtrip4 m1_5438_n3340#
+ m1_24338_n3340# m1_2792_4059# vtrip7 m1_2792_4059# m1_23582_n3340# m1_5438_n3340#
+ m1_4304_4059# vtrip4 vtrip6 m1_23960_4059# m1_20180_4059# avss m1_9596_4059# m1_17156_4059#
+ m1_23582_n3340# m1_12620_4059# m1_7706_n3340# m1_25472_4059# m1_5816_4059# m1_902_n3340#
+ m1_6950_n3340# m1_13376_4059# m1_22070_n3340# m1_9218_n3340# m1_2414_n3340# m1_9218_n3340#
+ m1_11486_n3340# m1_10352_4059# m1_17912_4059# m1_2414_n3340# m1_1280_4059# m1_24716_4059#
+ m1_10730_n3340# m1_6572_4059# m1_21692_4059# vtrip3 m1_9596_4059# m1_17912_4059#
+ m1_18290_n3340# m1_24716_4059# m1_25094_n3340# m1_2036_4059# vtrip6 m1_4682_n3340#
+ m1_20936_4059# m1_17156_4059# m1_8840_4059# m1_4682_n3340# m1_12620_4059# m1_3548_4059#
+ m1_25472_4059# sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2
Xsky130_fd_pr__nfet_g5v0d10v5_CD9S2Z_0 avss avss vtop ena_b sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
.ends

.subckt schmitt_trigger in out dvdd dvss
Xsky130_fd_pr__nfet_01v8_SCV3UK_1 m out dvss dvss m dvss dvss dvss in out m in sky130_fd_pr__nfet_01v8_SCV3UK
Xsky130_fd_pr__pfet_01v8_BZXTE7_0 dvdd dvdd out m out m in out dvdd dvdd m in dvdd
+ in m m in m out dvdd dvdd in m out m in dvdd dvdd sky130_fd_pr__pfet_01v8_BZXTE7
.ends

.subckt sky130_fd_pr__pfet_01v8_MA8JJJ a_18_n136# a_n33_95# w_n112_n198# a_n76_n136#
X0 a_18_n136# a_n33_95# a_n76_n136# w_n112_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_V6VPPZ a_n1842_n10916# a_n708_n10916# a_426_10484#
+ a_804_10484# a_n1464_n10916# a_n1972_n11046# a_1182_10484# a_n1086_n10916# a_1560_10484#
+ a_48_n10916# a_804_n10916# a_n330_10484# a_n708_10484# a_1560_n10916# a_48_10484#
+ a_426_n10916# a_n1086_10484# a_n1464_10484# a_1182_n10916# a_n1842_10484# a_n330_n10916#
X0 a_426_10484# a_426_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X1 a_n708_10484# a_n708_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X2 a_1560_10484# a_1560_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X3 a_n1086_10484# a_n1086_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X4 a_n1842_10484# a_n1842_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X5 a_n330_10484# a_n330_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X6 a_1182_10484# a_1182_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X7 a_48_10484# a_48_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X8 a_804_10484# a_804_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X9 a_n1464_10484# a_n1464_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
.ends

.subckt sky130_fd_pr__pfet_01v8_LAUYMQ w_n161_n200# a_n125_n100# a_66_n100# a_15_131#
+ a_n30_n100# a_n81_n197#
X0 a_n30_n100# a_n81_n197# a_n125_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.18
X1 a_66_n100# a_15_131# a_n30_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.18
.ends

.subckt sky130_fd_pr__pfet_01v8_C64SS5 a_287_n64# a_n187_n64# a_129_n64# w_n539_n164#
+ a_29_n161# a_n129_n161# a_187_n161# a_n29_n64# a_n287_n161# a_n503_n64# a_345_n161#
+ a_n345_n64# a_445_n64# a_n445_n161#
X0 a_129_n64# a_29_n161# a_n29_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n64# a_n287_n161# a_n345_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n345_n64# a_n445_n161# a_n503_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n29_n64# a_n129_n161# a_n187_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_287_n64# a_187_n161# a_129_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_445_n64# a_345_n161# a_287_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_2XUZHN a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_C68ZY6 a_208_n64# a_n108_n64# a_108_n161# w_n618_n164#
+ a_50_n64# a_n208_n161# a_266_n161# a_n424_n64# a_524_n64# a_n366_n161# a_424_n161#
+ a_n266_n64# a_366_n64# a_n524_n161# a_n50_n161# a_n582_n64#
X0 a_50_n64# a_n50_n161# a_n108_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n266_n64# a_n366_n161# a_n424_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n424_n64# a_n524_n161# a_n582_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n108_n64# a_n208_n161# a_n266_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_366_n64# a_266_n161# a_208_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_524_n64# a_424_n161# a_366_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X6 a_208_n64# a_108_n161# a_50_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_C6GQGA w_n154_n164# a_n118_n64# a_60_n64# a_n60_n161#
X0 a_60_n64# a_n60_n161# a_n118_n64# w_n154_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.6
.ends

.subckt sky130_fd_pr__pfet_01v8_9QCJ55 a_358_n64# a_n158_n64# a_158_n161# a_n358_n161#
+ a_n100_n161# w_n452_n164# a_100_n64# a_n416_n64#
X0 a_100_n64# a_n100_n161# a_n158_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 a_358_n64# a_158_n161# a_100_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2 a_n158_n64# a_n358_n161# a_n416_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_MLERZ7 a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt rc_osc dvdd out ena dvss
Xsky130_fd_pr__pfet_01v8_MA8JJJ_0 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_MA8JJJ
Xsky130_fd_pr__res_xhigh_po_1p41_V6VPPZ_0 vr m1_2270_n4# m1_23669_n1138# m1_23669_n1138#
+ m1_2270_752# dvss m1_23669_n1894# m1_2270_752# m1_23669_n1894# m1_2270_n760# m1_2270_n1516#
+ m1_23669_n382# m1_23669_374# in m1_23669_n382# m1_2270_n760# m1_23669_374# m1_23669_1130#
+ m1_2270_n1516# m1_23669_1130# m1_2270_n4# sky130_fd_pr__res_xhigh_po_1p41_V6VPPZ
Xsky130_fd_pr__pfet_01v8_LAUYMQ_0 dvdd dvdd vr ena_b out dvdd sky130_fd_pr__pfet_01v8_LAUYMQ
Xsky130_fd_pr__pfet_01v8_C64SS5_0 m dvdd dvdd dvdd in in in m in dvdd in m dvdd in
+ sky130_fd_pr__pfet_01v8_C64SS5
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 in dvdd dvdd ena sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_C68ZY6_0 out n n dvdd dvdd m n n out m n dvdd dvdd dvdd m
+ m sky130_fd_pr__pfet_01v8_C68ZY6
Xsky130_fd_pr__pfet_01v8_C6GQGA_0 dvdd dvdd ena_b ena sky130_fd_pr__pfet_01v8_C6GQGA
Xsky130_fd_pr__pfet_01v8_9QCJ55_0 m m n n n dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_9QCJ55
Xsky130_fd_pr__pfet_01v8_MLERZ7_0 vr ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_MLERZ7
X0 dvss dvss m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 m n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 dvss ena ena_b dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 out ena vr dvss sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X4 dvss dvss n dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 dvss in m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 n m dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 dvss dvss out dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X8 m in dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X9 vr dvss dvss dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X10 out n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_75J6LY a_n3403_n597# a_5977_n500# a_5177_n597#
+ a_29_n597# a_n2603_n500# a_5119_n500# a_n6893_n500# a_3461_n597# a_3403_n500# a_n6035_n500#
+ a_n2545_n597# w_n7093_n797# a_n1745_n500# a_4319_n597# a_n6835_n597# a_2545_n500#
+ a_2603_n597# a_n5177_n500# a_n1687_n597# a_n4261_n597# a_n887_n500# a_6835_n500#
+ a_n3461_n500# a_6035_n597# a_n5977_n597# a_n29_n500# a_n5119_n597# a_1687_n500#
+ a_1745_n597# a_n829_n597# a_4261_n500# a_887_n597# a_829_n500# a_n4319_n500#
X0 a_n6035_n500# a_n6835_n597# a_n6893_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1 a_3403_n500# a_2603_n597# a_2545_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_n29_n500# a_n829_n597# a_n887_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X3 a_n5177_n500# a_n5977_n597# a_n6035_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_2545_n500# a_1745_n597# a_1687_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_4261_n500# a_3461_n597# a_3403_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X6 a_n4319_n500# a_n5119_n597# a_n5177_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X7 a_829_n500# a_29_n597# a_n29_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X8 a_n2603_n500# a_n3403_n597# a_n3461_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X9 a_1687_n500# a_887_n597# a_829_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X10 a_6835_n500# a_6035_n597# a_5977_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X11 a_5119_n500# a_4319_n597# a_4261_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X12 a_n3461_n500# a_n4261_n597# a_n4319_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X13 a_n1745_n500# a_n2545_n597# a_n2603_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X14 a_5977_n500# a_5177_n597# a_5119_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X15 a_n887_n500# a_n1687_n597# a_n1745_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
.ends

.subckt ibias_gen ibias0 itest ibias1 ibg_200n vbg_1v2 isrc_sel ena ve avss avdd
Xsky130_fd_pr__nfet_g5v0d10v5_XZ4X25_0 isrc_sel_b ena_b isrc_sel avss ena_b vn1 avss
+ avss avss vn0 sky130_fd_pr__nfet_g5v0d10v5_XZ4X25
Xsky130_fd_pr__pfet_g5v0d10v5_Y9S9FP_0 avdd ena vp0 isrc_sel vp1 avdd avdd vp ena
+ avdd ena isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP
Xsky130_fd_pr__nfet_g5v0d10v5_62W3XE_0 avss isrc_sel isrc_sel_b ena_b ena avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_62W3XE
Xsky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1 vp0 vstart isrc_sel avss vn0 isrc_sel vbg_1v2
+ vn0 vn0 avss ibg_200n vn0 vbg_1v2 vp1 avss vbg_1v2 vstart isrc_sel_b vbg_1v2 vstart
+ vp vbg_1v2 avss vn0 vn1 vbg_1v2 vbg_1v2 vp vn0 vstart vbg_1v2 vstart ena vbg_1v2
+ vbg_1v2 sky130_fd_pr__nfet_g5v0d10v5_EC8RE7
Xsky130_fd_pr__pfet_g5v0d10v5_Y9J9EP_0 ena avdd avdd isrc_sel_b ena_b isrc_sel avdd
+ avdd sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP
Xsky130_fd_pr__nfet_g5v0d10v5_QZVU2P_1 avss vr ve avss avss vn0 avss vp0 avss ve avss
+ vn0 vn0 vn0 vr vn0 sky130_fd_pr__nfet_g5v0d10v5_QZVU2P
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_4165_119# m1_3409_119# m1_3409_119# m1_5299_7518#
+ m1_1519_7518# m1_385_119# m1_2653_119# m1_385_119# m1_2653_119# m1_6433_119# m1_1897_119#
+ avss m1_6055_7518# m1_3787_7518# m1_2275_7518# m1_1519_7518# m1_6055_7518# m1_4165_119#
+ m1_5299_7518# m1_763_7518# m1_4921_119# m1_763_7518# m1_7189_119# m1_4543_7518#
+ m1_1897_119# m1_7189_119# m1_3031_7518# m1_6811_7518# m1_4921_119# m1_5677_119#
+ m1_5677_119# m1_6811_7518# m1_3031_7518# m1_3787_7518# m1_1141_119# avss m1_4543_7518#
+ m1_1141_119# m1_6433_119# vr m1_2275_7518# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0 vn1 isrc_sel vp avdd vp1 vstart isrc_sel_b
+ ena_b avdd ibg_200n avdd isrc_sel ena_b avdd vp0 vp avdd isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_7JLQGA
Xsky130_fd_pr__nfet_g5v0d10v5_3DCHX4_0 avss avss vn1 avss avss avss avss avss vn1
+ avss avss avss vn1 avss avss avss vn1 vn1 avss vn1 vp1 avss avss avss avss vp1 avss
+ vn1 avss avss avss avss avss vn1 avss vp1 avss vp1 avss vn1 vn1 avss vn1 avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_3DCHX4
Xsky130_fd_pr__pfet_g5v0d10v5_75J6LY_0 vp0 avdd vp vp vp0 ibias1 avdd vp1 vp1 avdd
+ vp0 avdd avdd vp avdd avdd vp1 vn0 avdd avdd avdd avdd avdd avdd vp0 ibias0 vp0
+ itest vp vp avdd vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5_75J6LY
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5HVT2F a_1629_n430# a_4945_n65# a_n3287_n1257#
+ a_n3287_n892# a_3345_n162# a_4945_665# a_n3287_568# w_n5203_n1457# a_3345_n1257#
+ a_3287_1030# a_n1629_933# a_n5003_1030# a_3287_n1160# a_n29_n795# a_n4945_n527#
+ a_n1687_1030# a_3345_933# a_n4945_933# a_1687_n1257# a_4945_n430# a_1687_n527# a_n1629_568#
+ a_29_933# a_29_n527# a_3345_568# a_n4945_568# a_n5003_n1160# a_3345_n892# a_n3345_300#
+ a_n3345_n1160# a_n3345_n795# a_n1687_n65# a_n1629_n162# a_29_568# a_29_n1257# a_1629_n795#
+ a_n3287_n527# a_3287_300# a_n29_300# a_n1687_665# a_n29_1030# a_n1687_n1160# a_3287_n430#
+ a_n5003_n430# a_n1687_n430# a_n4945_n162# a_4945_n795# a_1687_n162# a_1629_300#
+ a_n5003_300# a_n1629_n892# a_1687_203# a_4945_300# a_n3287_203# a_1629_1030# a_n3345_1030#
+ a_3345_n527# a_n3345_n65# a_29_n162# a_n3345_665# a_n4945_n1257# a_n4945_n892# a_n29_n430#
+ a_3287_n65# a_n29_n65# a_n29_665# a_n3287_n162# a_3287_665# a_4945_n1160# a_3287_n795#
+ a_n5003_n795# a_1687_n892# a_n1629_203# a_4945_1030# a_n1629_n1257# a_1687_933#
+ a_n1687_n795# a_3345_203# a_n4945_203# a_n3287_933# a_n29_n1160# a_29_n892# a_1629_n1160#
+ a_n1629_n527# a_1629_n65# a_n5003_n65# a_1629_665# a_n5003_665# a_n3345_n430# a_n1687_300#
+ a_29_203# a_1687_568#
X0 a_n29_665# a_n1629_568# a_n1687_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n3345_n795# a_n4945_n892# a_n5003_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2 a_n29_300# a_n1629_203# a_n1687_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_4945_n430# a_3345_n527# a_3287_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X4 a_3287_n795# a_1687_n892# a_1629_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X5 a_n29_1030# a_n1629_933# a_n1687_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n1687_n795# a_n3287_n892# a_n3345_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n3345_665# a_n4945_568# a_n5003_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X8 a_n3345_300# a_n4945_203# a_n5003_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X9 a_n1687_n65# a_n3287_n162# a_n3345_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X10 a_n29_n1160# a_n1629_n1257# a_n1687_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_1629_665# a_29_568# a_n29_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X12 a_4945_n795# a_3345_n892# a_3287_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X13 a_n29_n430# a_n1629_n527# a_n1687_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_3287_665# a_1687_568# a_1629_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X15 a_1629_1030# a_29_933# a_n29_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_1629_300# a_29_203# a_n29_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X17 a_4945_665# a_3345_568# a_3287_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X18 a_3287_300# a_1687_203# a_1629_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X19 a_n29_n65# a_n1629_n162# a_n1687_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_n3345_1030# a_n4945_933# a_n5003_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X21 a_4945_300# a_3345_203# a_3287_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X22 a_3287_1030# a_1687_933# a_1629_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n3345_n65# a_n4945_n162# a_n5003_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X24 a_n1687_1030# a_n3287_933# a_n3345_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X25 a_n29_n795# a_n1629_n892# a_n1687_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X26 a_n3345_n1160# a_n4945_n1257# a_n5003_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X27 a_1629_n430# a_29_n527# a_n29_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X28 a_n1687_n1160# a_n3287_n1257# a_n3345_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X29 a_4945_n1160# a_3345_n1257# a_3287_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X30 a_1629_n65# a_29_n162# a_n29_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X31 a_n3345_n430# a_n4945_n527# a_n5003_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X32 a_4945_1030# a_3345_933# a_3287_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X33 a_n1687_665# a_n3287_568# a_n3345_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X34 a_3287_n65# a_1687_n162# a_1629_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 a_3287_n430# a_1687_n527# a_1629_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X36 a_1629_n1160# a_29_n1257# a_n29_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X37 a_n1687_n430# a_n3287_n527# a_n3345_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X38 a_n1687_300# a_n3287_203# a_n3345_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X39 a_4945_n65# a_3345_n162# a_3287_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X40 a_1629_n795# a_29_n892# a_n29_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X41 a_3287_n1160# a_1687_n1257# a_1629_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZV8547 a_3345_439# a_3287_527# a_1687_21# a_n4945_439#
+ a_n5003_n1563# a_1629_n1145# a_3345_n815# a_3287_n727# a_29_439# a_n5003_n727# a_n3345_n1563#
+ a_n4945_1275# a_n29_1363# a_4945_n309# a_3345_n397# a_n1687_n727# a_1687_1275# a_n1687_n1563#
+ a_n5003_527# a_1629_527# a_n4945_n1651# a_29_n1233# a_3287_n1145# a_n3345_109# a_29_1275#
+ a_4945_527# a_n1687_945# a_n3287_21# a_n29_109# a_3287_109# a_n3345_1363# a_29_21#
+ a_n5003_n1145# a_n1629_n1651# a_n1629_n815# a_1629_1363# a_n3287_1275# a_1687_857#
+ a_3287_n309# a_n29_n727# a_n5003_n309# a_n3345_n1145# a_n3287_857# a_n1629_n397#
+ a_n1687_n309# a_n1687_n1145# a_n5003_109# a_1629_109# a_n4945_n815# a_n4945_n1233#
+ a_n3287_n1651# a_4945_1363# a_n4945_21# a_4945_n1563# a_n3345_945# a_1687_n815#
+ a_3345_n1651# a_n1629_21# a_4945_109# a_n1687_527# a_n4945_n397# a_n3345_n727# a_n1629_857#
+ a_3345_1275# a_n29_n1563# a_1629_n727# a_1687_n1651# a_29_n815# a_n29_945# a_n1629_n1233#
+ a_1687_n397# a_3345_857# a_3287_945# a_n4945_857# a_3345_21# a_1629_n1563# a_1687_439#
+ a_n29_n309# a_29_n397# a_29_857# a_n3287_439# a_n3287_n815# a_3287_1363# a_n5003_1363#
+ a_4945_n727# a_n5137_n1785# a_n3287_n1233# a_n1687_1363# a_n5003_945# a_1629_945#
+ a_4945_n1145# a_29_n1651# a_3287_n1563# a_n3345_527# a_n3287_n397# a_3345_n1233#
+ a_4945_945# a_n1687_109# a_n1629_1275# a_n3345_n309# a_n1629_439# a_n29_n1145# a_1629_n309#
+ a_1687_n1233# a_n29_527#
X0 a_n1687_527# a_n3287_439# a_n3345_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_3287_n1563# a_1687_n1651# a_1629_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 a_3287_945# a_1687_857# a_1629_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_1629_109# a_29_21# a_n29_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_4945_945# a_3345_857# a_3287_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X5 a_3287_109# a_1687_21# a_1629_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_4945_n727# a_3345_n815# a_3287_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X7 a_4945_109# a_3345_21# a_3287_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X8 a_n29_527# a_n1629_439# a_n1687_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_n3345_n1145# a_n4945_n1233# a_n5003_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X10 a_n29_1363# a_n1629_1275# a_n1687_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_1629_n309# a_29_n397# a_n29_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X12 a_n1687_n1145# a_n3287_n1233# a_n3345_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X13 a_n3345_527# a_n4945_439# a_n5003_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X14 a_4945_n1145# a_3345_n1233# a_3287_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X15 a_n29_n1563# a_n1629_n1651# a_n1687_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_n3345_n309# a_n4945_n397# a_n5003_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X17 a_3287_n309# a_1687_n397# a_1629_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X18 a_n29_n727# a_n1629_n815# a_n1687_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X19 a_1629_n1145# a_29_n1233# a_n29_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_n1687_n309# a_n3287_n397# a_n3345_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n1687_945# a_n3287_857# a_n3345_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X22 a_1629_527# a_29_439# a_n29_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n1687_109# a_n3287_21# a_n3345_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X24 a_3287_n1145# a_1687_n1233# a_1629_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X25 a_1629_1363# a_29_1275# a_n29_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X26 a_3287_527# a_1687_439# a_1629_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X27 a_4945_527# a_3345_439# a_3287_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X28 a_4945_n309# a_3345_n397# a_3287_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X29 a_n3345_1363# a_n4945_1275# a_n5003_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X30 a_n29_945# a_n1629_857# a_n1687_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X31 a_3287_1363# a_1687_1275# a_1629_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X32 a_n29_109# a_n1629_21# a_n1687_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X33 a_n3345_n1563# a_n4945_n1651# a_n5003_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X34 a_n1687_1363# a_n3287_1275# a_n3345_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 a_1629_n727# a_29_n815# a_n29_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X36 a_n1687_n1563# a_n3287_n1651# a_n3345_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X37 a_4945_n1563# a_3345_n1651# a_3287_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X38 a_n3345_945# a_n4945_857# a_n5003_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X39 a_n3345_n727# a_n4945_n815# a_n5003_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X40 a_n3345_109# a_n4945_21# a_n5003_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X41 a_3287_n727# a_1687_n815# a_1629_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X42 a_n29_n1145# a_n1629_n1233# a_n1687_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X43 a_1629_n1563# a_29_n1651# a_n29_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X44 a_n1687_n727# a_n3287_n815# a_n3345_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X45 a_n29_n309# a_n1629_n397# a_n1687_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X46 a_4945_1363# a_3345_1275# a_3287_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X47 a_1629_945# a_29_857# a_n29_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5HV9F5 a_1629_118# a_n5003_118# a_1687_21# a_n29_n612#
+ a_n3287_n344# a_4945_118# a_29_386# a_n1687_483# a_n29_n247# a_n3345_n612# a_n1629_n709#
+ a_1629_n612# a_3345_n344# a_29_21# a_n3287_21# a_n3345_n247# a_n3345_483# w_n5203_n909#
+ a_n4945_n709# a_1629_n247# a_4945_n612# a_n1687_118# a_1687_n709# a_3287_483# a_n29_483#
+ a_29_n709# a_n4945_21# a_n1629_21# a_4945_n247# a_n1629_n344# a_n3287_n709# a_1629_483#
+ a_n5003_483# a_3345_21# a_1687_386# a_3287_n612# a_n5003_n612# a_n3345_118# a_4945_483#
+ a_n3287_386# a_n1687_n612# a_n4945_n344# a_n29_118# a_3287_n247# a_n5003_n247# a_1687_n344#
+ a_3287_118# a_n1687_n247# a_n1629_386# a_3345_n709# a_29_n344# a_3345_386# a_n4945_386#
X0 a_4945_n247# a_3345_n344# a_3287_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1 a_4945_n612# a_3345_n709# a_3287_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2 a_n29_118# a_n1629_21# a_n1687_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_n1687_483# a_n3287_386# a_n3345_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_n3345_118# a_n4945_21# a_n5003_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X5 a_n29_483# a_n1629_386# a_n1687_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n29_n612# a_n1629_n709# a_n1687_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n29_n247# a_n1629_n344# a_n1687_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X8 a_1629_118# a_29_21# a_n29_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_n3345_483# a_n4945_386# a_n5003_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X10 a_3287_118# a_1687_21# a_1629_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_4945_118# a_3345_21# a_3287_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X12 a_1629_483# a_29_386# a_n29_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X13 a_1629_n247# a_29_n344# a_n29_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_1629_n612# a_29_n709# a_n29_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X15 a_3287_483# a_1687_386# a_1629_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_n3345_n247# a_n4945_n344# a_n5003_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X17 a_n3345_n612# a_n4945_n709# a_n5003_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X18 a_4945_483# a_3345_386# a_3287_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X19 a_3287_n612# a_1687_n709# a_1629_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_3287_n247# a_1687_n344# a_1629_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n1687_n247# a_n3287_n344# a_n3345_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X22 a_n1687_n612# a_n3287_n709# a_n3345_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n1687_118# a_n3287_21# a_n3345_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt comparator ibias out ena vinn vinp avss vt avdd
Xsky130_fd_pr__pfet_g5v0d10v5_5H9LZ4_0 ena avdd ena vn vpp ena_b ena_b ibias ena avdd
+ vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4
Xsky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0 avdd vm vnn avdd avdd vpp avdd vpp avdd avdd
+ vnn n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5_3HV7M9
Xsky130_fd_pr__nfet_g5v0d10v5_T82T27_1 n0 vm vm avss vn avss avss avss vm vm vn avss
+ avss vn vn avss avss vn vm avss avss avss avss avss avss vt avss sky130_fd_pr__nfet_g5v0d10v5_T82T27
Xsky130_fd_pr__pfet_g5v0d10v5_5HVT2F_0 vnn avdd vnn vnn avdd avdd vnn avdd avdd avdd
+ vnn avdd avdd avdd avdd vpp avdd avdd vpp avdd vpp vnn vpp vpp avdd avdd avdd avdd
+ avdd avdd avdd vpp vnn vpp vpp vnn vnn avdd avdd vpp avdd vpp avdd avdd vpp avdd
+ avdd vpp vnn avdd vnn vpp avdd vnn vnn avdd avdd avdd vpp avdd avdd avdd avdd avdd
+ avdd avdd vnn avdd avdd avdd avdd vpp vnn avdd vnn vpp vpp avdd avdd vnn avdd vpp
+ vnn vnn vnn avdd vnn avdd avdd vpp vpp vpp sky130_fd_pr__pfet_g5v0d10v5_5HVT2F
Xsky130_fd_pr__nfet_g5v0d10v5_GG9S2Z_0 ena vm vn vn avss ena_b ena n0 avss avss ena_b
+ ibias avss ena_b avss ena_b sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z
Xsky130_fd_pr__nfet_g5v0d10v5_HZHY2Z_0 avss n1 n1 avss n1 avss n1 n1 out avss n0 avss
+ n1 n0 avss out n1 n1 out avss out n1 sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_ZV8547_0 avss vnn vinn avss vt vt avss vnn vinp vt vnn
+ avss vpp vt avss vt vinn vt vt vt avss vinp vnn vnn vinp vt vt vinn vpp vnn vnn
+ vinp vt vinp vinp vt vinn vinn vnn vpp vt vnn vinn vinp vt vt vt vt avss avss vinn
+ vt avss vt vnn vinn avss vinp vt vt avss vnn vinp avss vpp vt vinn vinp vpp vinp
+ vinn avss vnn avss avss vt vinn vpp vinp vinp vinn vinn vnn vt vt vt vinn vt vt
+ vt vt vinp vnn vnn vinn avss vt vt vinp vnn vinp vpp vt vinn vpp sky130_fd_pr__nfet_g5v0d10v5_ZV8547
Xsky130_fd_pr__pfet_g5v0d10v5_5HV9F5_0 vnn avdd vnn avdd vpp avdd vnn vpp avdd avdd
+ vpp vnn avdd vnn vpp avdd avdd avdd avdd vnn avdd vpp vnn avdd avdd vnn avdd vpp
+ avdd vpp vpp vnn avdd avdd vnn avdd avdd avdd avdd vpp vpp avdd avdd avdd avdd vnn
+ avdd vpp vpp avdd vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5HV9F5
Xsky130_fd_pr__pfet_g5v0d10v5_W8MWAU_0 out avdd avdd n1 n1 avdd n1 n1 avdd n1 out
+ n1 avdd n1 avdd n1 n0 out n1 out n0 avdd sky130_fd_pr__pfet_g5v0d10v5_W8MWAU
.ends

.subckt brownout_ana otrip_decoded[7] otrip_decoded[5] otrip_decoded[3] otrip_decoded[1]
+ vin_vunder vbg_1v2 ena ibg_200n itest isrc_sel vtrip_decoded[7] vtrip_decoded[6]
+ vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2] vtrip_decoded[0]
+ dcomp brout_filt osc_ena vunder outb comparator_1/vt otrip_decoded[4] dvdd comparator_0/vt
+ otrip_decoded[2] osc_ck outb_unbuf avdd vtrip_decoded[1] otrip_decoded[6] otrip_decoded[0]
+ avss vin_brout dvss
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_4_4/Y dvss dvss dvdd dvdd outb sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hvl__lsbufhv2lv_1_0 dcomp3v3 dvdd dvss dvss avdd avdd vl sky130_fd_sc_hvl__lsbufhv2lv_1
Xsky130_fd_sc_hvl__lsbufhv2lv_1_1 dcomp3v3uv dvdd dvss dvss avdd avdd sky130_fd_sc_hd__inv_4_2/A
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xrstring_mux_0 vin_brout ibias_gen_0/ena rstring_mux_0/otrip_decoded_avdd[7] rstring_mux_0/otrip_decoded_avdd[6]
+ rstring_mux_0/otrip_decoded_avdd[5] rstring_mux_0/otrip_decoded_avdd[4] rstring_mux_0/otrip_decoded_avdd[3]
+ rstring_mux_0/otrip_decoded_avdd[2] rstring_mux_0/otrip_decoded_avdd[1] rstring_mux_0/vtrip_decoded_avdd[7]
+ rstring_mux_0/vtrip_decoded_avdd[6] rstring_mux_0/vtrip_decoded_avdd[5] rstring_mux_0/vtrip_decoded_avdd[4]
+ rstring_mux_0/vtrip_decoded_avdd[3] rstring_mux_0/vtrip_decoded_avdd[2] rstring_mux_0/vtrip_decoded_avdd[1]
+ rstring_mux_0/vtrip_decoded_avdd[0] vin_vunder rstring_mux_0/vtop rstring_mux_0/otrip_decoded_avdd[0]
+ avdd avss rstring_mux
Xsky130_fd_sc_hd__inv_4_0 schmitt_trigger_0/out dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_0/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_1 sky130_fd_sc_hd__inv_4_2/Y dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_2 sky130_fd_sc_hd__inv_4_2/A dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_2/Y
+ sky130_fd_sc_hd__inv_4
Xschmitt_trigger_0 schmitt_trigger_0/in schmitt_trigger_0/out dvdd dvss schmitt_trigger
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] otrip_decoded[0] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] otrip_decoded[1] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] otrip_decoded[2] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] otrip_decoded[3] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2] otrip_decoded[4] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2] otrip_decoded[5] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3] otrip_decoded[6] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3] otrip_decoded[7] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4] vtrip_decoded[0] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4] vtrip_decoded[1] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5] vtrip_decoded[2] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5] vtrip_decoded[3] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6] vtrip_decoded[4] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6] vtrip_decoded[5] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7] vtrip_decoded[6] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7] vtrip_decoded[7] dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8] ena dvdd dvss dvss avdd avdd ibias_gen_0/ena
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8] isrc_sel dvdd dvss dvss avdd avdd ibias_gen_0/isrc_sel
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xrc_osc_0 dvdd osc_ck osc_ena dvss rc_osc
Xsky130_fd_sc_hd__inv_4_3 vl dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_4 outb_unbuf dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_4/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_n11325_2001# m1_n11325_2001# m1_n12081_2001#
+ m1_n10191_9400# m1_n13971_9400# m1_n14349_2001# m1_n12081_2001# vl m1_n12837_2001#
+ m1_n8301_2001# m1_n12837_2001# avss m1_n9435_9400# m1_n10947_9400# m1_n13215_9400#
+ m1_n13215_9400# m1_n8679_9400# m1_n10569_2001# m1_n9435_9400# m1_n13971_9400# m1_n10569_2001#
+ m1_n14727_9400# m1_n8301_2001# m1_n10947_9400# m1_n13593_2001# schmitt_trigger_0/in
+ m1_n11703_9400# m1_n8679_9400# m1_n9813_2001# m1_n9057_2001# m1_n9813_2001# m1_n7923_9400#
+ m1_n12459_9400# m1_n11703_9400# m1_n13593_2001# m1_n14727_9400# m1_n10191_9400#
+ m1_n14349_2001# m1_n9057_2001# m1_n7923_9400# m1_n12459_9400# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 schmitt_trigger_0/in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xibias_gen_0 ibias_gen_0/ibias0 itest ibias_gen_0/ibias1 ibg_200n vbg_1v2 ibias_gen_0/isrc_sel
+ ibias_gen_0/ena ibias_gen_0/ve avss avdd ibias_gen
Xsky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 avss avss ibias_gen_0/ve sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 m=1
Xcomparator_0 ibias_gen_0/ibias1 dcomp3v3uv ibias_gen_0/ena vin_vunder vbg_1v2 avss
+ comparator_0/vt avdd comparator
Xcomparator_1 ibias_gen_0/ibias0 dcomp3v3 ibias_gen_0/ena vin_brout vbg_1v2 avss comparator_1/vt
+ avdd comparator
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_4_0/Y dvss dvss dvdd dvdd brout_filt
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_4_1/Y dvss dvss dvdd dvdd vunder sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_4_3/Y dvss dvss dvdd dvdd dcomp sky130_fd_sc_hd__inv_16
.ends

.subckt sky130_ajc_ip__brownout avdd outb dvdd osc_ck dcomp vbg_1v2 otrip[2] otrip[1]
+ otrip[0] itest brout_filt vtrip[2] vtrip[1] vtrip[0] vin_brout ena force_ena_rc_osc
+ vin_vunder force_dis_rc_osc timed_out vunder force_short_oneshot isrc_sel ibg_200n
+ brownout_ana_0/comparator_1/vt brownout_ana_0/comparator_0/vt avss dvss
Xsky130_fd_pr__nfet_g5v0d10v5_PXF6AN_0 dvss dvss ena dvss dvss dvss dvss dvss dvss
+ dvss otrip[1] dvss dvss force_short_oneshot dvss dvss dvss dvss dvss force_dis_rc_osc
+ dvss otrip[2] force_ena_rc_osc dvss dvss dvss dvss otrip[0] isrc_sel dvss dvss dvss
+ dvss dvss sky130_fd_pr__nfet_g5v0d10v5_PXF6AN
Xbrownout_dig_0 dvdd brout_filt dcomp ena force_dis_rc_osc force_ena_rc_osc force_short_oneshot
+ osc_ck otrip[0] otrip[1] otrip[2] vtrip[0] vtrip[1] vtrip[2] brownout_dig_0/osc_ena
+ brownout_dig_0/otrip_decoded[0] brownout_dig_0/otrip_decoded[1] brownout_dig_0/otrip_decoded[3]
+ brownout_dig_0/otrip_decoded[4] brownout_dig_0/otrip_decoded[5] brownout_dig_0/otrip_decoded[6]
+ brownout_dig_0/otrip_decoded[7] brownout_dig_0/outb_unbuf timed_out brownout_dig_0/vtrip_decoded[0]
+ brownout_dig_0/vtrip_decoded[1] brownout_dig_0/vtrip_decoded[2] brownout_dig_0/vtrip_decoded[3]
+ brownout_dig_0/vtrip_decoded[4] brownout_dig_0/vtrip_decoded[5] brownout_dig_0/vtrip_decoded[6]
+ brownout_dig_0/vtrip_decoded[7] brownout_dig_0/otrip_decoded[2] dvss brownout_dig
Xsky130_fd_pr__nfet_g5v0d10v5_V6EN4F_0 dvss vin_vunder dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_V6EN4F
Xsky130_fd_pr__nfet_g5v0d10v5_XTZQRT_0 dvss dvss vtrip[1] dvss dvss dvss dvss dvss
+ dvss dvss vin_brout dvss dvss dvss dvss vbg_1v2 vtrip[2] dvss dvss dvss vtrip[0]
+ dvss sky130_fd_pr__nfet_g5v0d10v5_XTZQRT
Xbrownout_ana_0 brownout_dig_0/otrip_decoded[7] brownout_dig_0/otrip_decoded[5] brownout_dig_0/otrip_decoded[3]
+ brownout_dig_0/otrip_decoded[1] vin_vunder vbg_1v2 ena ibg_200n itest isrc_sel brownout_dig_0/vtrip_decoded[7]
+ brownout_dig_0/vtrip_decoded[6] brownout_dig_0/vtrip_decoded[5] brownout_dig_0/vtrip_decoded[4]
+ brownout_dig_0/vtrip_decoded[3] brownout_dig_0/vtrip_decoded[2] brownout_dig_0/vtrip_decoded[0]
+ dcomp brout_filt brownout_dig_0/osc_ena vunder outb brownout_ana_0/comparator_1/vt
+ brownout_dig_0/otrip_decoded[4] dvdd brownout_ana_0/comparator_0/vt brownout_dig_0/otrip_decoded[2]
+ osc_ck brownout_dig_0/outb_unbuf avdd brownout_dig_0/vtrip_decoded[1] brownout_dig_0/otrip_decoded[6]
+ brownout_dig_0/otrip_decoded[0] avss vin_brout dvss brownout_ana
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_W75H7K a_n4673_n1200# a_4873_n1200# a_2093_n1264#
+ a_n4099_n1264# w_n5131_n1497# a_4099_n1200# a_745_n1200# a_1577_n1264# a_803_n1264#
+ a_n745_n1264# a_n1003_n1264# a_n545_n1200# a_4157_n1264# a_n3583_n1264# a_3583_n1200#
+ a_1003_n1200# a_n3383_n1200# a_n2867_n1200# a_3641_n1264# a_n2293_n1264# a_2293_n1200#
+ a_n1577_n1200# a_n2093_n1200# a_n4931_n1200# a_2351_n1264# a_n1777_n1264# a_n4357_n1264#
+ a_1777_n1200# a_n29_n1200# a_n4157_n1200# a_1835_n1264# a_4357_n1200# a_n803_n1200#
+ a_4415_n1264# a_n3841_n1264# a_229_n1200# a_n3641_n1200# a_n229_n1264# a_3841_n1200#
+ a_1061_n1264# a_n3067_n1264# a_3067_n1200# a_3125_n1264# a_n2551_n1264# a_n2351_n1200#
+ a_2609_n1264# a_2551_n1200# a_n1835_n1200# a_n4615_n1264# a_4615_n1200# a_n4415_n1200#
+ a_1319_n1264# a_n1261_n1264# a_1261_n1200# a_n1061_n1200# a_3899_n1264# a_287_n1264#
+ a_n3325_n1264# a_n3125_n1200# a_n2809_n1264# a_3325_n1200# a_n2609_n1200# a_2809_n1200#
+ a_n2035_n1264# a_2035_n1200# a_n1519_n1264# a_1519_n1200# a_n1319_n1200# a_487_n1200#
+ a_n3899_n1200# a_4673_n1264# a_545_n1264# a_29_n1264# a_n487_n1264# a_n287_n1200#
+ a_3383_n1264# a_2867_n1264# a_n4873_n1264#
X0 a_3067_n1200# a_2867_n1264# a_2809_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X1 a_1777_n1200# a_1577_n1264# a_1519_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X2 a_2809_n1200# a_2609_n1264# a_2551_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X3 a_n4157_n1200# a_n4357_n1264# a_n4415_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X4 a_1519_n1200# a_1319_n1264# a_1261_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X5 a_4873_n1200# a_4673_n1264# a_4615_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=1.74 ps=12.29 w=12 l=1
X6 a_3583_n1200# a_3383_n1264# a_3325_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X7 a_4615_n1200# a_4415_n1264# a_4357_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X8 a_n2867_n1200# a_n3067_n1264# a_n3125_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X9 a_487_n1200# a_287_n1264# a_229_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X10 a_2293_n1200# a_2093_n1264# a_2035_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X11 a_3325_n1200# a_3125_n1264# a_3067_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X12 a_n287_n1200# a_n487_n1264# a_n545_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X13 a_n2609_n1200# a_n2809_n1264# a_n2867_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X14 a_n1577_n1200# a_n1777_n1264# a_n1835_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X15 a_n29_n1200# a_n229_n1264# a_n287_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X16 a_n4673_n1200# a_n4873_n1264# a_n4931_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=3.48 ps=24.58 w=12 l=1
X17 a_n1319_n1200# a_n1519_n1264# a_n1577_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X18 a_2035_n1200# a_1835_n1264# a_1777_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X19 a_n4415_n1200# a_n4615_n1264# a_n4673_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X20 a_n3383_n1200# a_n3583_n1264# a_n3641_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X21 a_n3125_n1200# a_n3325_n1264# a_n3383_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X22 a_3841_n1200# a_3641_n1264# a_3583_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X23 a_n2093_n1200# a_n2293_n1264# a_n2351_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X24 a_745_n1200# a_545_n1264# a_487_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X25 a_2551_n1200# a_2351_n1264# a_2293_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X26 a_n1835_n1200# a_n2035_n1264# a_n2093_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X27 a_1261_n1200# a_1061_n1264# a_1003_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X28 a_n545_n1200# a_n745_n1264# a_n803_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X29 a_229_n1200# a_29_n1264# a_n29_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X30 a_4099_n1200# a_3899_n1264# a_3841_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X31 a_n3641_n1200# a_n3841_n1264# a_n3899_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X32 a_n2351_n1200# a_n2551_n1264# a_n2609_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X33 a_1003_n1200# a_803_n1264# a_745_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X34 a_n3899_n1200# a_n4099_n1264# a_n4157_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X35 a_n1061_n1200# a_n1261_n1264# a_n1319_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X36 a_4357_n1200# a_4157_n1264# a_4099_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X37 a_n803_n1200# a_n1003_n1264# a_n1061_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CVG6CD a_50_n400# w_n308_n697# a_n50_n464# a_n108_n400#
X0 a_50_n400# a_n50_n464# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WKXP7K a_n4673_n1200# a_4873_n1200# a_4931_n1264#
+ a_2093_n1264# a_n4099_n1264# a_4099_n1200# a_745_n1200# a_1577_n1264# a_803_n1264#
+ a_n745_n1264# a_n1003_n1264# a_n545_n1200# a_4157_n1264# a_n3583_n1264# a_3583_n1200#
+ a_1003_n1200# a_n3383_n1200# a_n2867_n1200# a_3641_n1264# a_n2293_n1264# a_2293_n1200#
+ a_n1577_n1200# a_n2093_n1200# a_n4931_n1200# a_2351_n1264# a_n1777_n1264# a_n4357_n1264#
+ a_1777_n1200# a_n29_n1200# a_n4157_n1200# a_1835_n1264# a_4357_n1200# a_n803_n1200#
+ a_4415_n1264# a_n3841_n1264# a_229_n1200# a_n3641_n1200# a_n229_n1264# a_3841_n1200#
+ a_1061_n1264# a_n3067_n1264# a_3067_n1200# a_3125_n1264# a_n2551_n1264# a_n2351_n1200#
+ a_2609_n1264# a_n5131_n1264# w_n5389_n1497# a_5131_n1200# a_2551_n1200# a_n1835_n1200#
+ a_n4615_n1264# a_4615_n1200# a_n4415_n1200# a_1319_n1264# a_n1261_n1264# a_1261_n1200#
+ a_n1061_n1200# a_3899_n1264# a_287_n1264# a_n3325_n1264# a_n3125_n1200# a_n2809_n1264#
+ a_3325_n1200# a_n2609_n1200# a_2809_n1200# a_n2035_n1264# a_2035_n1200# a_n1519_n1264#
+ a_1519_n1200# a_n1319_n1200# a_487_n1200# a_n3899_n1200# a_4673_n1264# a_545_n1264#
+ a_29_n1264# a_n487_n1264# a_n287_n1200# a_3383_n1264# a_n5189_n1200# a_2867_n1264#
+ a_n4873_n1264#
X0 a_3067_n1200# a_2867_n1264# a_2809_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X1 a_1777_n1200# a_1577_n1264# a_1519_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X2 a_2809_n1200# a_2609_n1264# a_2551_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X3 a_n4157_n1200# a_n4357_n1264# a_n4415_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X4 a_1519_n1200# a_1319_n1264# a_1261_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X5 a_4873_n1200# a_4673_n1264# a_4615_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X6 a_3583_n1200# a_3383_n1264# a_3325_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X7 a_4615_n1200# a_4415_n1264# a_4357_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X8 a_n2867_n1200# a_n3067_n1264# a_n3125_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X9 a_487_n1200# a_287_n1264# a_229_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X10 a_2293_n1200# a_2093_n1264# a_2035_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X11 a_3325_n1200# a_3125_n1264# a_3067_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X12 a_n287_n1200# a_n487_n1264# a_n545_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X13 a_n2609_n1200# a_n2809_n1264# a_n2867_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X14 a_n1577_n1200# a_n1777_n1264# a_n1835_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X15 a_n29_n1200# a_n229_n1264# a_n287_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X16 a_n4673_n1200# a_n4873_n1264# a_n4931_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X17 a_n1319_n1200# a_n1519_n1264# a_n1577_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X18 a_2035_n1200# a_1835_n1264# a_1777_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X19 a_5131_n1200# a_4931_n1264# a_4873_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=1.74 ps=12.29 w=12 l=1
X20 a_n4415_n1200# a_n4615_n1264# a_n4673_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X21 a_n3383_n1200# a_n3583_n1264# a_n3641_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X22 a_n3125_n1200# a_n3325_n1264# a_n3383_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X23 a_3841_n1200# a_3641_n1264# a_3583_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X24 a_n2093_n1200# a_n2293_n1264# a_n2351_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X25 a_745_n1200# a_545_n1264# a_487_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X26 a_2551_n1200# a_2351_n1264# a_2293_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X27 a_n1835_n1200# a_n2035_n1264# a_n2093_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X28 a_n4931_n1200# a_n5131_n1264# a_n5189_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=3.48 ps=24.58 w=12 l=1
X29 a_1261_n1200# a_1061_n1264# a_1003_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X30 a_n545_n1200# a_n745_n1264# a_n803_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X31 a_229_n1200# a_29_n1264# a_n29_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X32 a_4099_n1200# a_3899_n1264# a_3841_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X33 a_n3641_n1200# a_n3841_n1264# a_n3899_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X34 a_n2351_n1200# a_n2551_n1264# a_n2609_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X35 a_1003_n1200# a_803_n1264# a_745_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X36 a_n3899_n1200# a_n4099_n1264# a_n4157_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X37 a_n1061_n1200# a_n1261_n1264# a_n1319_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X38 a_4357_n1200# a_4157_n1264# a_4099_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X39 a_n803_n1200# a_n1003_n1264# a_n1061_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_6H2JYD a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CTEUHA a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HQ4STX w_n358_n597# a_n158_n300# a_n100_n364#
+ a_100_n300#
X0 a_100_n300# a_n100_n364# a_n158_n300# w_n358_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J a_1519_n450# a_n803_n450# a_n2093_n450#
+ a_n2551_n505# a_1261_n450# a_29_n505# a_n1777_n505# a_n3067_n505# a_n1319_n450#
+ a_n287_n450# a_n1061_n450# a_2867_n505# a_n745_n505# a_2809_n450# a_803_n505# a_n2035_n505#
+ a_745_n450# a_n3383_n450# a_2551_n450# a_3125_n505# a_1835_n505# a_3067_n450# a_1777_n450#
+ a_n2609_n450# a_n229_n505# a_n1003_n505# a_n2351_n450# a_287_n505# a_2093_n505#
+ a_229_n450# a_n1577_n450# a_n3325_n505# a_2035_n450# a_1319_n505# a_n545_n450# a_1061_n505#
+ a_n2293_n505# a_n3517_n672# a_1003_n450# a_n1519_n505# a_n2867_n450# a_n487_n505#
+ a_3325_n450# a_n1261_n505# a_2609_n505# a_n29_n450# a_545_n505# a_487_n450# a_2351_n505#
+ a_2293_n450# a_n1835_n450# a_n3125_n450# a_1577_n505# a_n2809_n505#
X0 a_n2351_n450# a_n2551_n505# a_n2609_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X1 a_n2093_n450# a_n2293_n505# a_n2351_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X2 a_229_n450# a_29_n505# a_n29_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X3 a_n29_n450# a_n229_n505# a_n287_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X4 a_3067_n450# a_2867_n505# a_2809_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X5 a_n1319_n450# a_n1519_n505# a_n1577_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X6 a_n545_n450# a_n745_n505# a_n803_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X7 a_2551_n450# a_2351_n505# a_2293_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X8 a_n3125_n450# a_n3325_n505# a_n3383_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=1
X9 a_n287_n450# a_n487_n505# a_n545_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X10 a_2293_n450# a_2093_n505# a_2035_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X11 a_n2867_n450# a_n3067_n505# a_n3125_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X12 a_n803_n450# a_n1003_n505# a_n1061_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X13 a_n1577_n450# a_n1777_n505# a_n1835_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X14 a_1519_n450# a_1319_n505# a_1261_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X15 a_n1061_n450# a_n1261_n505# a_n1319_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X16 a_3325_n450# a_3125_n505# a_3067_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=1
X17 a_1003_n450# a_803_n505# a_745_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X18 a_745_n450# a_545_n505# a_487_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X19 a_487_n450# a_287_n505# a_229_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X20 a_2035_n450# a_1835_n505# a_1777_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X21 a_n2609_n450# a_n2809_n505# a_n2867_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X22 a_1777_n450# a_1577_n505# a_1519_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X23 a_1261_n450# a_1061_n505# a_1003_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X24 a_n1835_n450# a_n2035_n505# a_n2093_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X25 a_2809_n450# a_2609_n505# a_2551_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_USXRNR a_1448_n255# a_1190_n255# a_358_n200#
+ a_n1648_n255# a_n1706_n200# a_100_n200# a_n674_n200# a_n616_n255# a_n1390_n255#
+ a_674_n255# a_1132_n200# a_n158_n200# a_158_n255# a_616_n200# a_n874_n255# a_n932_n200#
+ a_1648_n200# a_932_n255# a_1390_n200# a_n1448_n200# a_n358_n255# a_n416_n200# a_n1190_n200#
+ a_n1132_n255# a_874_n200# a_416_n255# a_n100_n255# a_n1840_n422#
X0 a_1648_n200# a_1448_n255# a_1390_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X1 a_1132_n200# a_932_n255# a_874_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_874_n200# a_674_n255# a_616_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1390_n200# a_1190_n255# a_1132_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_100_n200# a_n100_n255# a_n158_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n416_n200# a_n616_n255# a_n674_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n158_n200# a_n358_n255# a_n416_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n1448_n200# a_n1648_n255# a_n1706_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X8 a_n1190_n200# a_n1390_n255# a_n1448_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n674_n200# a_n874_n255# a_n932_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n932_n200# a_n1132_n255# a_n1190_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_358_n200# a_158_n255# a_100_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_616_n200# a_416_n255# a_358_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AUMBFF a_n2035_n2564# a_n1519_n2564# a_2035_n2500#
+ a_n1319_n2500# a_1519_n2500# a_n3899_n2500# a_487_n2500# a_545_n2564# a_29_n2564#
+ a_n487_n2564# a_n287_n2500# a_3383_n2564# a_2867_n2564# a_2093_n2564# a_n4099_n2564#
+ a_745_n2500# a_1577_n2564# a_803_n2564# a_n1003_n2564# w_n4615_n2797# a_4099_n2500#
+ a_n545_n2500# a_4157_n2564# a_n745_n2564# a_n3583_n2564# a_1003_n2500# a_n3383_n2500#
+ a_3583_n2500# a_n2867_n2500# a_3641_n2564# a_n2293_n2564# a_2293_n2500# a_n2093_n2500#
+ a_n1777_n2564# a_1777_n2500# a_n29_n2500# a_n1577_n2500# a_n4157_n2500# a_2351_n2564#
+ a_n4357_n2564# a_4357_n2500# a_1835_n2564# a_229_n2500# a_n803_n2500# a_n229_n2564#
+ a_n3841_n2564# a_3841_n2500# a_n3641_n2500# a_1061_n2564# a_n3067_n2564# a_3067_n2500#
+ a_3125_n2564# a_n2551_n2564# a_n2351_n2500# a_2609_n2564# a_2551_n2500# a_n1835_n2500#
+ a_n4415_n2500# a_1319_n2564# a_n1261_n2564# a_1261_n2500# a_n1061_n2500# a_3899_n2564#
+ a_n3125_n2500# a_287_n2564# a_n2809_n2564# a_n3325_n2564# a_3325_n2500# a_n2609_n2500#
+ a_2809_n2500#
X0 a_3067_n2500# a_2867_n2564# a_2809_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X1 a_2809_n2500# a_2609_n2564# a_2551_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X2 a_1777_n2500# a_1577_n2564# a_1519_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X3 a_n4157_n2500# a_n4357_n2564# a_n4415_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=7.25 ps=50.58 w=25 l=1
X4 a_1519_n2500# a_1319_n2564# a_1261_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X5 a_3583_n2500# a_3383_n2564# a_3325_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X6 a_n2867_n2500# a_n3067_n2564# a_n3125_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X7 a_487_n2500# a_287_n2564# a_229_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X8 a_2293_n2500# a_2093_n2564# a_2035_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X9 a_3325_n2500# a_3125_n2564# a_3067_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X10 a_n287_n2500# a_n487_n2564# a_n545_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X11 a_n2609_n2500# a_n2809_n2564# a_n2867_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X12 a_n1577_n2500# a_n1777_n2564# a_n1835_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X13 a_n29_n2500# a_n229_n2564# a_n287_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X14 a_2035_n2500# a_1835_n2564# a_1777_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X15 a_n1319_n2500# a_n1519_n2564# a_n1577_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X16 a_n3383_n2500# a_n3583_n2564# a_n3641_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X17 a_3841_n2500# a_3641_n2564# a_3583_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X18 a_n3125_n2500# a_n3325_n2564# a_n3383_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X19 a_n2093_n2500# a_n2293_n2564# a_n2351_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X20 a_745_n2500# a_545_n2564# a_487_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X21 a_n1835_n2500# a_n2035_n2564# a_n2093_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X22 a_2551_n2500# a_2351_n2564# a_2293_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X23 a_1261_n2500# a_1061_n2564# a_1003_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X24 a_n545_n2500# a_n745_n2564# a_n803_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X25 a_229_n2500# a_29_n2564# a_n29_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X26 a_4099_n2500# a_3899_n2564# a_3841_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X27 a_n3641_n2500# a_n3841_n2564# a_n3899_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X28 a_n2351_n2500# a_n2551_n2564# a_n2609_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X29 a_1003_n2500# a_803_n2564# a_745_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X30 a_n3899_n2500# a_n4099_n2564# a_n4157_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X31 a_n1061_n2500# a_n1261_n2564# a_n1319_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X32 a_n803_n2500# a_n1003_n2564# a_n1061_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X33 a_4357_n2500# a_4157_n2564# a_4099_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=7.25 pd=50.58 as=3.625 ps=25.29 w=25 l=1
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_25PWK4 a_n148_n148# a_n46_n46#
X0 a_n148_n148# a_n46_n46# sky130_fd_pr__diode_pw2nd_05v5 perim=1.84e+06 area=2.116e+11
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QL2RRT a_29_n664# a_n1777_n664# a_n2351_n600#
+ a_n745_n664# a_229_n600# a_n1577_n600# a_2867_n664# a_2035_n600# a_803_n664# a_n2035_n664#
+ a_n545_n600# a_3125_n664# a_1835_n664# a_1003_n600# a_n229_n664# w_n3583_n897# a_287_n664#
+ a_n1003_n664# a_n2867_n600# a_3325_n600# a_2093_n664# a_n3325_n664# a_n29_n600#
+ a_487_n600# a_1319_n664# a_2293_n600# a_n3125_n600# a_n2293_n664# a_n1835_n600#
+ a_1061_n664# a_n803_n600# a_1519_n600# a_n2093_n600# a_n1519_n664# a_1261_n600#
+ a_n487_n664# a_n1261_n664# a_2609_n664# a_545_n664# a_n1319_n600# a_n287_n600# a_n1061_n600#
+ a_2351_n664# a_2809_n600# a_1577_n664# a_745_n600# a_n3383_n600# a_n2809_n664# a_2551_n600#
+ a_n2551_n664# a_3067_n600# a_1777_n600# a_n2609_n600# a_n3067_n664#
X0 a_n1835_n600# a_n2035_n664# a_n2093_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_2809_n600# a_2609_n664# a_2551_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2351_n600# a_n2551_n664# a_n2609_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_n2093_n600# a_n2293_n664# a_n2351_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_229_n600# a_29_n664# a_n29_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_n29_n600# a_n229_n664# a_n287_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_3067_n600# a_2867_n664# a_2809_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_n1319_n600# a_n1519_n664# a_n1577_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n545_n600# a_n745_n664# a_n803_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X9 a_2551_n600# a_2351_n664# a_2293_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n3125_n600# a_n3325_n664# a_n3383_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X11 a_n287_n600# a_n487_n664# a_n545_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_2293_n600# a_2093_n664# a_2035_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n2867_n600# a_n3067_n664# a_n3125_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n803_n600# a_n1003_n664# a_n1061_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_n1577_n600# a_n1777_n664# a_n1835_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_1519_n600# a_1319_n664# a_1261_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_n1061_n600# a_n1261_n664# a_n1319_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X18 a_3325_n600# a_3125_n664# a_3067_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X19 a_1003_n600# a_803_n664# a_745_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_487_n600# a_287_n664# a_229_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_745_n600# a_545_n664# a_487_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_2035_n600# a_1835_n664# a_1777_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_n2609_n600# a_n2809_n664# a_n2867_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1777_n600# a_1577_n664# a_1519_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_1261_n600# a_1061_n664# a_1003_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_U4BBJH a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QTY6KC a_287_n464# a_n1003_n464# a_487_n400#
+ a_n29_n400# a_1319_n464# w_n1777_n697# a_1061_n464# a_1519_n400# a_n803_n400# a_n1519_n464#
+ a_1261_n400# a_n487_n464# a_n1261_n464# a_n1319_n400# a_545_n464# a_n287_n400# a_n1061_n400#
+ a_745_n400# a_29_n464# a_n745_n464# a_229_n400# a_n1577_n400# a_803_n464# a_n545_n400#
+ a_1003_n400# a_n229_n464#
X0 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_n545_n400# a_n745_n464# a_n803_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n287_n400# a_n487_n464# a_n545_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_1519_n400# a_1319_n464# a_1261_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X5 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_1003_n400# a_803_n464# a_745_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_487_n400# a_287_n464# a_229_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_745_n400# a_545_n464# a_487_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_1261_n400# a_1061_n464# a_1003_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n29_n400# a_n229_n464# a_n287_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_229_n400# a_29_n464# a_n29_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z a_1519_n450# a_n803_n450# a_n2093_n450#
+ a_n2551_n505# a_1261_n450# a_29_n505# a_n1777_n505# a_n3067_n505# a_n1319_n450#
+ a_3641_n505# a_3583_n450# a_n4033_n672# a_n287_n450# a_n1061_n450# a_2867_n505#
+ a_n745_n505# a_2809_n450# a_803_n505# a_n2035_n505# a_745_n450# a_n3383_n450# a_n3841_n505#
+ a_2551_n450# a_3125_n505# a_1835_n505# a_3067_n450# a_1777_n450# a_n2609_n450# a_n229_n505#
+ a_n1003_n505# a_n2351_n450# a_287_n505# a_2093_n505# a_229_n450# a_n1577_n450# a_n3325_n505#
+ a_2035_n450# a_3841_n450# a_1319_n505# a_n545_n450# a_n3899_n450# a_1061_n505# a_n2293_n505#
+ a_1003_n450# a_n3641_n450# a_3383_n505# a_n1519_n505# a_n2867_n450# a_n487_n505#
+ a_3325_n450# a_n1261_n505# a_2609_n505# a_n29_n450# a_545_n505# a_487_n450# a_2351_n505#
+ a_n3583_n505# a_2293_n450# a_n1835_n450# a_n3125_n450# a_1577_n505# a_n2809_n505#
X0 a_n2351_n450# a_n2551_n505# a_n2609_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X1 a_n2093_n450# a_n2293_n505# a_n2351_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X2 a_229_n450# a_29_n505# a_n29_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X3 a_n29_n450# a_n229_n505# a_n287_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X4 a_3067_n450# a_2867_n505# a_2809_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X5 a_n1319_n450# a_n1519_n505# a_n1577_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X6 a_n545_n450# a_n745_n505# a_n803_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X7 a_2551_n450# a_2351_n505# a_2293_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X8 a_n3125_n450# a_n3325_n505# a_n3383_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X9 a_n287_n450# a_n487_n505# a_n545_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X10 a_2293_n450# a_2093_n505# a_2035_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X11 a_n2867_n450# a_n3067_n505# a_n3125_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X12 a_n803_n450# a_n1003_n505# a_n1061_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X13 a_n1577_n450# a_n1777_n505# a_n1835_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X14 a_n3641_n450# a_n3841_n505# a_n3899_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=1
X15 a_n3383_n450# a_n3583_n505# a_n3641_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X16 a_1519_n450# a_1319_n505# a_1261_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X17 a_n1061_n450# a_n1261_n505# a_n1319_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X18 a_3325_n450# a_3125_n505# a_3067_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X19 a_1003_n450# a_803_n505# a_745_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X20 a_745_n450# a_545_n505# a_487_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X21 a_487_n450# a_287_n505# a_229_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X22 a_2035_n450# a_1835_n505# a_1777_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X23 a_n2609_n450# a_n2809_n505# a_n2867_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X24 a_1777_n450# a_1577_n505# a_1519_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X25 a_3841_n450# a_3641_n505# a_3583_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=1
X26 a_3583_n450# a_3383_n505# a_3325_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X27 a_1261_n450# a_1061_n505# a_1003_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X28 a_n1835_n450# a_n2035_n505# a_n2093_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X29 a_2809_n450# a_2609_n505# a_2551_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QTY6H6 a_1261_n200# a_n487_n264# a_n1261_n264#
+ a_n1319_n200# a_545_n264# a_n287_n200# a_n1061_n200# a_745_n200# a_29_n264# a_229_n200#
+ a_n745_n264# a_n1577_n200# a_803_n264# a_n545_n200# a_1003_n200# a_n229_n264# a_n1003_n264#
+ a_287_n264# a_487_n200# a_n29_n200# a_1319_n264# a_1061_n264# w_n1777_n497# a_n803_n200#
+ a_1519_n200# a_n1519_n264#
X0 a_745_n200# a_545_n264# a_487_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1003_n200# a_803_n264# a_745_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_487_n200# a_287_n264# a_229_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1261_n200# a_1061_n264# a_1003_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n29_n200# a_n229_n264# a_n287_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_229_n200# a_29_n264# a_n29_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n1319_n200# a_n1519_n264# a_n1577_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X7 a_n545_n200# a_n745_n264# a_n803_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n803_n200# a_n1003_n264# a_n1061_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n287_n200# a_n487_n264# a_n545_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_1519_n200# a_1319_n264# a_1261_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X11 a_n1061_n200# a_n1261_n264# a_n1319_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_U73S5M a_229_n1000# a_n803_n1000# a_545_n1055#
+ a_29_n1055# a_n487_n1055# a_n4549_n1222# a_n3641_n1000# a_3841_n1000# a_3067_n1000#
+ a_3383_n1055# a_2867_n1055# a_2551_n1000# a_n2351_n1000# a_n1835_n1000# a_n4415_n1000#
+ a_2093_n1055# a_n4099_n1055# a_1577_n1055# a_803_n1055# a_n745_n1055# a_n1003_n1055#
+ a_n1061_n1000# a_4157_n1055# a_n3583_n1055# a_1261_n1000# a_n3125_n1000# a_3641_n1055#
+ a_3325_n1000# a_2809_n1000# a_n2609_n1000# a_n2293_n1055# a_n1777_n1055# a_2035_n1000#
+ a_2351_n1055# a_n4357_n1055# a_1519_n1000# a_n1319_n1000# a_n3899_n1000# a_1835_n1055#
+ a_487_n1000# a_n229_n1055# a_n3841_n1055# a_n287_n1000# a_1061_n1055# a_n3067_n1055#
+ a_3125_n1055# a_n2551_n1055# a_2609_n1055# a_1319_n1055# a_n1261_n1055# a_4099_n1000#
+ a_745_n1000# a_3899_n1055# a_1003_n1000# a_n545_n1000# a_287_n1055# a_n2809_n1055#
+ a_n3325_n1055# a_3583_n1000# a_n3383_n1000# a_n2867_n1000# a_n2035_n1055# a_n2093_n1000#
+ a_n1519_n1055# a_2293_n1000# a_n1577_n1000# a_4357_n1000# a_1777_n1000# a_n29_n1000#
+ a_n4157_n1000#
X0 a_3067_n1000# a_2867_n1055# a_2809_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X1 a_n1319_n1000# a_n1519_n1055# a_n1577_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X2 a_n545_n1000# a_n745_n1055# a_n803_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X3 a_2293_n1000# a_2093_n1055# a_2035_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X4 a_2551_n1000# a_2351_n1055# a_2293_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X5 a_n3125_n1000# a_n3325_n1055# a_n3383_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X6 a_n2867_n1000# a_n3067_n1055# a_n3125_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X7 a_n803_n1000# a_n1003_n1055# a_n1061_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X8 a_n287_n1000# a_n487_n1055# a_n545_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X9 a_n3641_n1000# a_n3841_n1055# a_n3899_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X10 a_n1577_n1000# a_n1777_n1055# a_n1835_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X11 a_1519_n1000# a_1319_n1055# a_1261_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X12 a_n3383_n1000# a_n3583_n1055# a_n3641_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X13 a_3325_n1000# a_3125_n1055# a_3067_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X14 a_n1061_n1000# a_n1261_n1055# a_n1319_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X15 a_745_n1000# a_545_n1055# a_487_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X16 a_1003_n1000# a_803_n1055# a_745_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X17 a_487_n1000# a_287_n1055# a_229_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X18 a_2035_n1000# a_1835_n1055# a_1777_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X19 a_4099_n1000# a_3899_n1055# a_3841_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X20 a_n2609_n1000# a_n2809_n1055# a_n2867_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X21 a_1777_n1000# a_1577_n1055# a_1519_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X22 a_3841_n1000# a_3641_n1055# a_3583_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X23 a_1261_n1000# a_1061_n1055# a_1003_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X24 a_3583_n1000# a_3383_n1055# a_3325_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X25 a_n4157_n1000# a_n4357_n1055# a_n4415_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X26 a_n3899_n1000# a_n4099_n1055# a_n4157_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X27 a_n1835_n1000# a_n2035_n1055# a_n2093_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X28 a_2809_n1000# a_2609_n1055# a_2551_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X29 a_n2351_n1000# a_n2551_n1055# a_n2609_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X30 a_4357_n1000# a_4157_n1055# a_4099_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X31 a_n2093_n1000# a_n2293_n1055# a_n2351_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X32 a_n29_n1000# a_n229_n1055# a_n287_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X33 a_229_n1000# a_29_n1055# a_n29_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PP2RNK a_29_n964# a_n2351_n900# a_229_n900# a_2867_n964#
+ a_n745_n964# a_n1577_n900# a_2035_n900# a_803_n964# a_n2035_n964# a_n545_n900# w_n3325_n1197#
+ a_1835_n964# a_1003_n900# a_n229_n964# a_n1003_n964# a_287_n964# a_n2867_n900# a_2093_n964#
+ a_487_n900# a_n29_n900# a_2293_n900# a_n3125_n900# a_1319_n964# a_n1835_n900# a_1061_n964#
+ a_n2293_n964# a_n803_n900# a_1519_n900# a_n2093_n900# a_n1519_n964# a_1261_n900#
+ a_n487_n964# a_n1261_n964# a_2609_n964# a_n1319_n900# a_545_n964# a_n287_n900# a_2351_n964#
+ a_n1061_n900# a_1577_n964# a_2809_n900# a_745_n900# a_n2809_n964# a_2551_n900# a_n2551_n964#
+ a_3067_n900# a_1777_n900# a_n2609_n900# a_n1777_n964# a_n3067_n964#
X0 a_n2609_n900# a_n2809_n964# a_n2867_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1 a_1261_n900# a_1061_n964# a_1003_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X2 a_n1835_n900# a_n2035_n964# a_n2093_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X3 a_2809_n900# a_2609_n964# a_2551_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X4 a_n2351_n900# a_n2551_n964# a_n2609_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 a_n2093_n900# a_n2293_n964# a_n2351_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 a_n29_n900# a_n229_n964# a_n287_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X7 a_229_n900# a_29_n964# a_n29_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 a_3067_n900# a_2867_n964# a_2809_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X9 a_n1319_n900# a_n1519_n964# a_n1577_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 a_2551_n900# a_2351_n964# a_2293_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X11 a_n545_n900# a_n745_n964# a_n803_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 a_n287_n900# a_n487_n964# a_n545_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X13 a_2293_n900# a_2093_n964# a_2035_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X14 a_n2867_n900# a_n3067_n964# a_n3125_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X15 a_n803_n900# a_n1003_n964# a_n1061_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X16 a_n1577_n900# a_n1777_n964# a_n1835_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 a_1519_n900# a_1319_n964# a_1261_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X18 a_n1061_n900# a_n1261_n964# a_n1319_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X19 a_1003_n900# a_803_n964# a_745_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X20 a_745_n900# a_545_n964# a_487_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X21 a_487_n900# a_287_n964# a_229_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X22 a_1777_n900# a_1577_n964# a_1519_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X23 a_2035_n900# a_1835_n964# a_1777_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_79TVLH a_3067_n300# a_1777_n300# a_n2609_n300#
+ a_1061_n355# a_n2293_n355# a_n2351_n300# a_229_n300# a_n1577_n300# a_n1519_n355#
+ a_2035_n300# a_n487_n355# a_n545_n300# a_n1261_n355# a_2609_n355# a_545_n355# a_n3517_n522#
+ a_2351_n355# a_1003_n300# a_1577_n355# a_n2867_n300# a_n2809_n355# a_3325_n300#
+ a_n2551_n355# a_487_n300# a_n29_n300# a_n3067_n355# a_29_n355# a_n1777_n355# a_2293_n300#
+ a_n1835_n300# a_n3125_n300# a_n745_n355# a_2867_n355# a_1519_n300# a_n803_n300#
+ a_n2093_n300# a_803_n355# a_n2035_n355# a_1261_n300# a_n1319_n300# a_3125_n355#
+ a_1835_n355# a_n287_n300# a_n229_n355# a_n1061_n300# a_287_n355# a_n1003_n355# a_2809_n300#
+ a_745_n300# a_2093_n355# a_n3383_n300# a_n3325_n355# a_2551_n300# a_1319_n355#
X0 a_2809_n300# a_2609_n355# a_2551_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1 a_n2351_n300# a_n2551_n355# a_n2609_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X2 a_n2093_n300# a_n2293_n355# a_n2351_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3 a_n29_n300# a_n229_n355# a_n287_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X4 a_229_n300# a_29_n355# a_n29_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X5 a_3067_n300# a_2867_n355# a_2809_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 a_n1319_n300# a_n1519_n355# a_n1577_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_n545_n300# a_n745_n355# a_n803_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X8 a_2293_n300# a_2093_n355# a_2035_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X9 a_2551_n300# a_2351_n355# a_2293_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X10 a_n3125_n300# a_n3325_n355# a_n3383_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X11 a_n2867_n300# a_n3067_n355# a_n3125_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X12 a_n803_n300# a_n1003_n355# a_n1061_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_n287_n300# a_n487_n355# a_n545_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X14 a_n1577_n300# a_n1777_n355# a_n1835_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X15 a_1519_n300# a_1319_n355# a_1261_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 a_3325_n300# a_3125_n355# a_3067_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X17 a_n1061_n300# a_n1261_n355# a_n1319_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X18 a_745_n300# a_545_n355# a_487_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X19 a_1003_n300# a_803_n355# a_745_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X20 a_487_n300# a_287_n355# a_229_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X21 a_2035_n300# a_1835_n355# a_1777_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 a_n2609_n300# a_n2809_n355# a_n2867_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X23 a_1777_n300# a_1577_n355# a_1519_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_1261_n300# a_1061_n355# a_1003_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X25 a_n1835_n300# a_n2035_n355# a_n2093_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2B7385 a_1261_n800# a_n1319_n800# a_1835_n855#
+ a_n287_n800# a_n229_n855# a_n1061_n800# a_287_n855# a_n1003_n855# a_2093_n855# a_745_n800#
+ a_1319_n855# a_1777_n800# a_n2293_n855# a_n2351_n800# a_1061_n855# a_229_n800# a_2035_n800#
+ a_n1577_n800# a_n1519_n855# a_n487_n855# a_n1261_n855# a_n545_n800# a_545_n855#
+ a_1003_n800# a_1577_n855# a_n2485_n1022# a_n29_n800# a_487_n800# a_2293_n800# a_29_n855#
+ a_n1777_n855# a_n1835_n800# a_n745_n855# a_n803_n800# a_1519_n800# a_n2093_n800#
+ a_803_n855# a_n2035_n855#
X0 a_n1577_n800# a_n1777_n855# a_n1835_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X1 a_1519_n800# a_1319_n855# a_1261_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2 a_n1061_n800# a_n1261_n855# a_n1319_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X3 a_1003_n800# a_803_n855# a_745_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X4 a_745_n800# a_545_n855# a_487_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X5 a_487_n800# a_287_n855# a_229_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X6 a_1777_n800# a_1577_n855# a_1519_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X7 a_2035_n800# a_1835_n855# a_1777_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X8 a_1261_n800# a_1061_n855# a_1003_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X9 a_n1835_n800# a_n2035_n855# a_n2093_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X10 a_n2093_n800# a_n2293_n855# a_n2351_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X11 a_n29_n800# a_n229_n855# a_n287_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X12 a_229_n800# a_29_n855# a_n29_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X13 a_n1319_n800# a_n1519_n855# a_n1577_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X14 a_n545_n800# a_n745_n855# a_n803_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X15 a_n287_n800# a_n487_n855# a_n545_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X16 a_2293_n800# a_2093_n855# a_2035_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X17 a_n803_n800# a_n1003_n855# a_n1061_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NT3TPY a_n287_n255# a_n345_n200# a_345_n255#
+ a_n445_n255# a_129_n200# a_n503_n200# a_287_n200# a_445_n200# a_n637_n422# a_n29_n200#
+ a_29_n255# a_n187_n200# a_n129_n255# a_187_n255#
X0 a_n187_n200# a_n287_n255# a_n345_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n255# a_129_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n255# a_n503_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_129_n200# a_29_n255# a_n29_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n255# a_287_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n29_n200# a_n129_n255# a_n187_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR a_n2093_n200# a_803_n255# a_n2035_n255#
+ a_n3841_n255# a_n5131_n255# a_1261_n200# a_n4357_n255# a_3583_n200# a_n1319_n200#
+ a_n4415_n200# a_4931_n255# a_3125_n255# a_1835_n255# a_n287_n200# a_n229_n255# a_4099_n200#
+ a_n1061_n200# a_287_n255# a_n1003_n255# a_2809_n200# a_745_n200# a_n3383_n200# a_2093_n255#
+ a_n3325_n255# a_2551_n200# a_3067_n200# a_4415_n255# a_1319_n255# a_4873_n200# a_1777_n200#
+ a_n2609_n200# a_n2293_n255# a_1061_n255# a_n5323_n422# a_n2351_n200# a_229_n200#
+ a_3383_n255# a_n1577_n200# a_n4673_n200# a_n1519_n255# a_n4615_n255# a_5131_n200#
+ a_3841_n200# a_2035_n200# a_n487_n255# a_n545_n200# a_n3899_n200# a_n5189_n200#
+ a_n1261_n255# a_4357_n200# a_2609_n255# a_545_n255# a_n3583_n255# a_n3641_n200#
+ a_2351_n255# a_1003_n200# a_n4099_n255# a_n4157_n200# a_4673_n255# a_1577_n255#
+ a_3325_n200# a_n2867_n200# a_n2809_n255# a_3899_n255# a_n2551_n255# a_487_n200#
+ a_n29_n200# a_n3067_n255# a_2293_n200# a_29_n255# a_n1777_n255# a_n4873_n255# a_n1835_n200#
+ a_n3125_n200# a_n4931_n200# a_3641_n255# a_4157_n255# a_n745_n255# a_n803_n200#
+ a_2867_n255# a_4615_n200# a_1519_n200#
X0 a_487_n200# a_287_n255# a_229_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_2035_n200# a_1835_n255# a_1777_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_4099_n200# a_3899_n255# a_3841_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n2609_n200# a_n2809_n255# a_n2867_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_1777_n200# a_1577_n255# a_1519_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_3841_n200# a_3641_n255# a_3583_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n4415_n200# a_n4615_n255# a_n4673_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_1261_n200# a_1061_n255# a_1003_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_3583_n200# a_3383_n255# a_3325_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n4157_n200# a_n4357_n255# a_n4415_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n3899_n200# a_n4099_n255# a_n4157_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1835_n200# a_n2035_n255# a_n2093_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_n4673_n200# a_n4873_n255# a_n4931_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_2809_n200# a_2609_n255# a_2551_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_n2351_n200# a_n2551_n255# a_n2609_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_4357_n200# a_4157_n255# a_4099_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_4615_n200# a_4415_n255# a_4357_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_n2093_n200# a_n2293_n255# a_n2351_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_n29_n200# a_n229_n255# a_n287_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_229_n200# a_29_n255# a_n29_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_3067_n200# a_2867_n255# a_2809_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X21 a_5131_n200# a_4931_n255# a_4873_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X22 a_4873_n200# a_4673_n255# a_4615_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X24 a_n545_n200# a_n745_n255# a_n803_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X25 a_2293_n200# a_2093_n255# a_2035_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 a_2551_n200# a_2351_n255# a_2293_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X27 a_n4931_n200# a_n5131_n255# a_n5189_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X28 a_n3125_n200# a_n3325_n255# a_n3383_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 a_n2867_n200# a_n3067_n255# a_n3125_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X31 a_n287_n200# a_n487_n255# a_n545_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X32 a_n3641_n200# a_n3841_n255# a_n3899_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_n1577_n200# a_n1777_n255# a_n1835_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 a_1519_n200# a_1319_n255# a_1261_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X35 a_n3383_n200# a_n3583_n255# a_n3641_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 a_3325_n200# a_3125_n255# a_3067_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X38 a_745_n200# a_545_n255# a_487_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X39 a_1003_n200# a_803_n255# a_745_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WK95DB a_n819_n450# a_n345_n450# a_29_n505# a_n129_n505#
+ a_187_n505# a_129_n450# a_n503_n450# a_n287_n505# a_345_n505# a_287_n450# a_n661_n450#
+ a_n445_n505# a_503_n505# a_445_n450# a_n603_n505# a_661_n505# a_603_n450# a_n761_n505#
+ a_761_n450# a_n953_n672# a_n29_n450# a_n187_n450#
X0 a_n345_n450# a_n445_n505# a_n503_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X1 a_129_n450# a_29_n505# a_n29_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X2 a_445_n450# a_345_n505# a_287_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X3 a_n503_n450# a_n603_n505# a_n661_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X4 a_n29_n450# a_n129_n505# a_n187_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X5 a_603_n450# a_503_n505# a_445_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X6 a_n661_n450# a_n761_n505# a_n819_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.5
X7 a_n187_n450# a_n287_n505# a_n345_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X8 a_761_n450# a_661_n505# a_603_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.5
X9 a_287_n450# a_187_n505# a_129_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3QL9S5 a_n50_n497# a_50_n400# w_n308_n697# a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PGZBW9 a_1061_n655# a_n2293_n655# a_n2351_n600#
+ a_229_n600# a_n1577_n600# a_n1519_n655# a_2035_n600# a_n487_n655# a_n1261_n655#
+ a_n545_n600# a_2609_n655# a_545_n655# a_2351_n655# a_n3517_n822# a_1003_n600# a_1577_n655#
+ a_n2867_n600# a_n2809_n655# a_3325_n600# a_n2551_n655# a_n29_n600# a_487_n600# a_n1777_n655#
+ a_n3067_n655# a_2293_n600# a_n3125_n600# a_29_n655# a_n1835_n600# a_2867_n655# a_n745_n655#
+ a_n803_n600# a_1519_n600# a_n2093_n600# a_803_n655# a_n2035_n655# a_1261_n600# a_3125_n655#
+ a_n1319_n600# a_1835_n655# a_n287_n600# a_n1061_n600# a_n229_n655# a_n1003_n655#
+ a_287_n655# a_2809_n600# a_2093_n655# a_745_n600# a_n3383_n600# a_n3325_n655# a_2551_n600#
+ a_3067_n600# a_1777_n600# a_n2609_n600# a_1319_n655#
X0 a_2809_n600# a_2609_n655# a_2551_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n655# a_n2609_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n655# a_n2351_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_229_n600# a_29_n655# a_n29_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_n29_n600# a_n229_n655# a_n287_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n655# a_2809_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n655# a_n1577_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n655# a_2293_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n655# a_n3383_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X9 a_n545_n600# a_n745_n655# a_n803_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n655# a_n545_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n655# a_2035_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n655# a_n3125_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n655# a_n1061_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n1577_n600# a_n1777_n655# a_n1835_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_1519_n600# a_1319_n655# a_1261_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_n1061_n600# a_n1261_n655# a_n1319_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_3325_n600# a_3125_n655# a_3067_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X18 a_1003_n600# a_803_n655# a_745_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_745_n600# a_545_n655# a_487_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_487_n600# a_287_n655# a_229_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_2035_n600# a_1835_n655# a_1777_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_n2609_n600# a_n2809_n655# a_n2867_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_1777_n600# a_1577_n655# a_1519_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1261_n600# a_1061_n655# a_1003_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_n1835_n600# a_n2035_n655# a_n2093_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD a_761_n400# a_503_n464# a_n29_n400# a_n603_n464#
+ a_661_n464# a_n187_n400# a_n761_n464# a_n819_n400# a_n345_n400# a_129_n400# a_n503_n400#
+ w_n1019_n697# a_287_n400# a_n661_n400# a_29_n464# a_n129_n464# a_187_n464# a_445_n400#
+ a_n287_n464# a_345_n464# a_603_n400# a_n445_n464#
X0 a_n503_n400# a_n603_n464# a_n661_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n464# a_n187_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n464# a_445_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n661_n400# a_n761_n464# a_n819_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n187_n400# a_n287_n464# a_n345_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_761_n400# a_661_n464# a_603_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_287_n400# a_187_n464# a_129_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n345_n400# a_n445_n464# a_n503_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_129_n400# a_29_n464# a_n29_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_445_n400# a_345_n464# a_287_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QSKB8C a_287_n464# a_n1003_n464# a_n2867_n400#
+ a_n4157_n400# a_2093_n464# a_3325_n400# a_n3325_n464# a_487_n400# a_n29_n400# a_4415_n464#
+ a_1319_n464# a_2293_n400# a_n1835_n400# a_n3125_n400# a_n2293_n464# a_n4931_n400#
+ a_1061_n464# a_1519_n400# a_n803_n400# a_3383_n464# a_4615_n400# a_n2093_n400# a_n1519_n464#
+ a_n4615_n464# a_1261_n400# a_n487_n464# a_n1261_n464# w_n5131_n697# a_n1319_n400#
+ a_2609_n464# a_545_n464# a_3583_n400# a_n287_n400# a_n4415_n400# a_n3583_n464# a_4099_n400#
+ a_n1061_n400# a_2351_n464# a_n4099_n464# a_2809_n400# a_4673_n464# a_1577_n464#
+ a_745_n400# a_n3383_n400# a_n2809_n464# a_2551_n400# a_3899_n464# a_n2551_n464#
+ a_4873_n400# a_3067_n400# a_1777_n400# a_n2609_n400# a_n3067_n464# a_3641_n464#
+ a_29_n464# a_n1777_n464# a_n4873_n464# a_n2351_n400# a_4157_n464# a_n745_n464# a_229_n400#
+ a_n1577_n400# a_n4673_n400# a_2867_n464# a_2035_n400# a_803_n464# a_n2035_n464#
+ a_3841_n400# a_n3841_n464# a_4357_n400# a_n545_n400# a_n3899_n400# a_3125_n464#
+ a_n4357_n464# a_1835_n464# a_1003_n400# a_n3641_n400# a_n229_n464#
X0 a_3067_n400# a_2867_n464# a_2809_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_4873_n400# a_4673_n464# a_4615_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n545_n400# a_n745_n464# a_n803_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_2293_n400# a_2093_n464# a_2035_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_2551_n400# a_2351_n464# a_2293_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n3125_n400# a_n3325_n464# a_n3383_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n2867_n400# a_n3067_n464# a_n3125_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_n287_n400# a_n487_n464# a_n545_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n3641_n400# a_n3841_n464# a_n3899_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_n1577_n400# a_n1777_n464# a_n1835_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_1519_n400# a_1319_n464# a_1261_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_n3383_n400# a_n3583_n464# a_n3641_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_3325_n400# a_3125_n464# a_3067_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_1003_n400# a_803_n464# a_745_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_487_n400# a_287_n464# a_229_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_745_n400# a_545_n464# a_487_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_2035_n400# a_1835_n464# a_1777_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_4099_n400# a_3899_n464# a_3841_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_n2609_n400# a_n2809_n464# a_n2867_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X22 a_1777_n400# a_1577_n464# a_1519_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X23 a_3841_n400# a_3641_n464# a_3583_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X24 a_n4415_n400# a_n4615_n464# a_n4673_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 a_1261_n400# a_1061_n464# a_1003_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X26 a_3583_n400# a_3383_n464# a_3325_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X27 a_n4157_n400# a_n4357_n464# a_n4415_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X28 a_n3899_n400# a_n4099_n464# a_n4157_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X29 a_n1835_n400# a_n2035_n464# a_n2093_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X30 a_n4673_n400# a_n4873_n464# a_n4931_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X31 a_2809_n400# a_2609_n464# a_2551_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X32 a_n2351_n400# a_n2551_n464# a_n2609_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X33 a_4357_n400# a_4157_n464# a_4099_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X34 a_4615_n400# a_4415_n464# a_4357_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X35 a_n2093_n400# a_n2293_n464# a_n2351_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X36 a_n29_n400# a_n229_n464# a_n287_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X37 a_229_n400# a_29_n464# a_n29_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QRKB8C a_287_n464# a_n1003_n464# a_n2867_n400#
+ a_n4157_n400# a_2093_n464# a_3325_n400# a_n3325_n464# a_487_n400# a_n29_n400# a_4415_n464#
+ a_1319_n464# a_2293_n400# a_n1835_n400# a_n3125_n400# a_n2293_n464# a_1061_n464#
+ w_n4873_n697# a_1519_n400# a_n803_n400# a_3383_n464# a_4615_n400# a_n2093_n400#
+ a_n1519_n464# a_n4615_n464# a_1261_n400# a_n487_n464# a_n1261_n464# a_n1319_n400#
+ a_2609_n464# a_545_n464# a_3583_n400# a_n287_n400# a_n4415_n400# a_n3583_n464# a_4099_n400#
+ a_n1061_n400# a_2351_n464# a_n4099_n464# a_2809_n400# a_1577_n464# a_745_n400# a_n3383_n400#
+ a_n2809_n464# a_2551_n400# a_3899_n464# a_n2551_n464# a_3067_n400# a_1777_n400#
+ a_n2609_n400# a_n3067_n464# a_3641_n464# a_29_n464# a_n1777_n464# a_n2351_n400#
+ a_4157_n464# a_n745_n464# a_229_n400# a_n1577_n400# a_n4673_n400# a_2867_n464# a_2035_n400#
+ a_803_n464# a_n2035_n464# a_3841_n400# a_n3841_n464# a_4357_n400# a_n545_n400# a_n3899_n400#
+ a_3125_n464# a_n4357_n464# a_1835_n464# a_1003_n400# a_n3641_n400# a_n229_n464#
X0 a_3067_n400# a_2867_n464# a_2809_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n545_n400# a_n745_n464# a_n803_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_2293_n400# a_2093_n464# a_2035_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_2551_n400# a_2351_n464# a_2293_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_n3125_n400# a_n3325_n464# a_n3383_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n2867_n400# a_n3067_n464# a_n3125_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n287_n400# a_n487_n464# a_n545_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_n3641_n400# a_n3841_n464# a_n3899_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n1577_n400# a_n1777_n464# a_n1835_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_1519_n400# a_1319_n464# a_1261_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_n3383_n400# a_n3583_n464# a_n3641_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_3325_n400# a_3125_n464# a_3067_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_1003_n400# a_803_n464# a_745_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_487_n400# a_287_n464# a_229_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_745_n400# a_545_n464# a_487_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_2035_n400# a_1835_n464# a_1777_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_4099_n400# a_3899_n464# a_3841_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_n2609_n400# a_n2809_n464# a_n2867_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_1777_n400# a_1577_n464# a_1519_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X22 a_3841_n400# a_3641_n464# a_3583_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X23 a_n4415_n400# a_n4615_n464# a_n4673_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X24 a_1261_n400# a_1061_n464# a_1003_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 a_3583_n400# a_3383_n464# a_3325_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X26 a_n4157_n400# a_n4357_n464# a_n4415_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X27 a_n3899_n400# a_n4099_n464# a_n4157_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X28 a_n1835_n400# a_n2035_n464# a_n2093_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X29 a_2809_n400# a_2609_n464# a_2551_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X30 a_n2351_n400# a_n2551_n464# a_n2609_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X31 a_4357_n400# a_4157_n464# a_4099_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X32 a_4615_n400# a_4415_n464# a_4357_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X33 a_n2093_n400# a_n2293_n464# a_n2351_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X34 a_n29_n400# a_n229_n464# a_n287_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X35 a_229_n400# a_29_n464# a_n29_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_Z5XS7R c1_6184_n8000# c1_n8876_n8000# m3_6144_n8040#
+ c1_160_n8000# m3_n2892_n8040# m3_n8916_n8040# c1_3172_n8000# c1_n5864_n8000# m3_3132_n8040#
+ m3_n5904_n8040# m3_120_n8040# c1_n2852_n8000#
X0 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X1 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X2 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X3 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X4 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X5 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X6 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X7 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X8 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X9 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X10 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X11 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X12 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X13 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X14 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X15 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X16 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X17 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X18 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X19 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X20 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X21 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X22 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X23 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X24 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X25 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X26 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X27 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X28 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X29 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X30 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X31 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X33 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X35 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_EVM3FM a_29_n964# a_n129_n964# a_187_n964# a_445_n900#
+ a_n287_n964# a_345_n964# a_603_n900# a_n445_n964# a_761_n900# a_503_n964# a_n29_n900#
+ a_n603_n964# a_661_n964# a_n187_n900# a_n761_n964# a_n819_n900# a_n345_n900# a_129_n900#
+ a_n503_n900# w_n1019_n1197# a_n661_n900# a_287_n900#
X0 a_n187_n900# a_n287_n964# a_n345_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X1 a_761_n900# a_661_n964# a_603_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=0.5
X2 a_287_n900# a_187_n964# a_129_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X3 a_n345_n900# a_n445_n964# a_n503_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X4 a_129_n900# a_29_n964# a_n29_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X5 a_445_n900# a_345_n964# a_287_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X6 a_n503_n900# a_n603_n964# a_n661_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X7 a_n29_n900# a_n129_n964# a_n187_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X8 a_603_n900# a_503_n964# a_445_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X9 a_n661_n900# a_n761_n964# a_n819_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN a_n2093_n200# a_803_n255# a_n2035_n255#
+ a_n3841_n255# a_1261_n200# a_n4357_n255# a_3583_n200# a_n1319_n200# a_n4415_n200#
+ a_3125_n255# a_1835_n255# a_n287_n200# a_n229_n255# a_4099_n200# a_n1061_n200# a_287_n255#
+ a_n1003_n255# a_2809_n200# a_745_n200# a_n3383_n200# a_2093_n255# a_n3325_n255#
+ a_2551_n200# a_3067_n200# a_4415_n255# a_1319_n255# a_4873_n200# a_1777_n200# a_n2609_n200#
+ a_n2293_n255# a_1061_n255# a_n2351_n200# a_229_n200# a_3383_n255# a_n1577_n200#
+ a_n4673_n200# a_n1519_n255# a_n4615_n255# a_3841_n200# a_2035_n200# a_n487_n255#
+ a_n545_n200# a_n3899_n200# a_n1261_n255# a_4357_n200# a_2609_n255# a_545_n255# a_n3583_n255#
+ a_n3641_n200# a_2351_n255# a_1003_n200# a_n4099_n255# a_n4157_n200# a_4673_n255#
+ a_1577_n255# a_3325_n200# a_n2867_n200# a_n2809_n255# a_3899_n255# a_n2551_n255#
+ a_487_n200# a_n29_n200# a_n3067_n255# a_2293_n200# a_29_n255# a_n1777_n255# a_n4873_n255#
+ a_n1835_n200# a_n3125_n200# a_n4931_n200# a_3641_n255# a_4157_n255# a_n745_n255#
+ a_n803_n200# a_2867_n255# a_4615_n200# a_1519_n200# a_n5065_n422#
X0 a_487_n200# a_287_n255# a_229_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_2035_n200# a_1835_n255# a_1777_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_4099_n200# a_3899_n255# a_3841_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n2609_n200# a_n2809_n255# a_n2867_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_1777_n200# a_1577_n255# a_1519_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_3841_n200# a_3641_n255# a_3583_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n4415_n200# a_n4615_n255# a_n4673_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_1261_n200# a_1061_n255# a_1003_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_3583_n200# a_3383_n255# a_3325_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n4157_n200# a_n4357_n255# a_n4415_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n3899_n200# a_n4099_n255# a_n4157_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1835_n200# a_n2035_n255# a_n2093_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_n4673_n200# a_n4873_n255# a_n4931_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X13 a_2809_n200# a_2609_n255# a_2551_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_n2351_n200# a_n2551_n255# a_n2609_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_4357_n200# a_4157_n255# a_4099_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_4615_n200# a_4415_n255# a_4357_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_n2093_n200# a_n2293_n255# a_n2351_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_n29_n200# a_n229_n255# a_n287_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_229_n200# a_29_n255# a_n29_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_3067_n200# a_2867_n255# a_2809_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X21 a_4873_n200# a_4673_n255# a_4615_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X22 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 a_n545_n200# a_n745_n255# a_n803_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X24 a_2293_n200# a_2093_n255# a_2035_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X25 a_2551_n200# a_2351_n255# a_2293_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 a_n3125_n200# a_n3325_n255# a_n3383_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X27 a_n2867_n200# a_n3067_n255# a_n3125_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X28 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 a_n287_n200# a_n487_n255# a_n545_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 a_n3641_n200# a_n3841_n255# a_n3899_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X31 a_n1577_n200# a_n1777_n255# a_n1835_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X32 a_1519_n200# a_1319_n255# a_1261_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_n3383_n200# a_n3583_n255# a_n3641_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 a_3325_n200# a_3125_n255# a_3067_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X35 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 a_745_n200# a_545_n255# a_487_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 a_1003_n200# a_803_n255# a_745_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Q46EE6 a_1261_n200# a_n487_n264# a_n1261_n264#
+ w_n2035_n497# a_n1319_n200# a_545_n264# a_n287_n200# a_n1061_n200# a_1577_n264#
+ a_745_n200# a_1777_n200# a_n1777_n264# a_29_n264# a_229_n200# a_n745_n264# a_n1577_n200#
+ a_803_n264# a_n545_n200# a_1003_n200# a_n229_n264# a_n1003_n264# a_287_n264# a_487_n200#
+ a_n29_n200# a_1319_n264# a_n1835_n200# a_1061_n264# a_n803_n200# a_1519_n200# a_n1519_n264#
X0 a_745_n200# a_545_n264# a_487_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1003_n200# a_803_n264# a_745_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_487_n200# a_287_n264# a_229_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1777_n200# a_1577_n264# a_1519_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X4 a_1261_n200# a_1061_n264# a_1003_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n29_n200# a_n229_n264# a_n287_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_229_n200# a_29_n264# a_n29_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n1319_n200# a_n1519_n264# a_n1577_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n545_n200# a_n745_n264# a_n803_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n803_n200# a_n1003_n264# a_n1061_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n287_n200# a_n487_n264# a_n545_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1577_n200# a_n1777_n264# a_n1835_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X12 a_1519_n200# a_1319_n264# a_1261_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_n1061_n200# a_n1261_n264# a_n1319_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UGZTXE a_1061_n655# a_n2293_n655# a_n2351_n600#
+ a_229_n600# a_n1577_n600# a_3383_n655# a_n1519_n655# a_2035_n600# a_n487_n655# a_n1261_n655#
+ a_n545_n600# a_2609_n655# a_545_n655# a_2351_n655# a_n3583_n655# a_1003_n600# a_n3641_n600#
+ a_1577_n655# a_n2867_n600# a_n2809_n655# a_3325_n600# a_n2551_n655# a_n29_n600#
+ a_487_n600# a_n1777_n655# a_n3067_n655# a_2293_n600# a_n3125_n600# a_29_n655# a_n1835_n600#
+ a_2867_n655# a_n745_n655# a_n803_n600# a_1519_n600# a_n2093_n600# a_803_n655# a_n2035_n655#
+ a_n3775_n822# a_1261_n600# a_3125_n655# a_3583_n600# a_n1319_n600# a_1835_n655#
+ a_n287_n600# a_n1061_n600# a_n229_n655# a_n1003_n655# a_287_n655# a_2809_n600# a_2093_n655#
+ a_745_n600# a_n3383_n600# a_n3325_n655# a_2551_n600# a_3067_n600# a_1777_n600# a_n2609_n600#
+ a_1319_n655#
X0 a_2809_n600# a_2609_n655# a_2551_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n655# a_n2609_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n655# a_n2351_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_229_n600# a_29_n655# a_n29_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_n29_n600# a_n229_n655# a_n287_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n655# a_2809_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n655# a_n1577_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n655# a_2293_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n655# a_n3383_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X9 a_n545_n600# a_n745_n655# a_n803_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n655# a_n545_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n655# a_2035_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n655# a_n3125_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n655# a_n1061_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n3383_n600# a_n3583_n655# a_n3641_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X15 a_n1577_n600# a_n1777_n655# a_n1835_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_1519_n600# a_1319_n655# a_1261_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_n1061_n600# a_n1261_n655# a_n1319_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X18 a_3325_n600# a_3125_n655# a_3067_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_1003_n600# a_803_n655# a_745_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_745_n600# a_545_n655# a_487_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_487_n600# a_287_n655# a_229_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_2035_n600# a_1835_n655# a_1777_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_n2609_n600# a_n2809_n655# a_n2867_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1777_n600# a_1577_n655# a_1519_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_3583_n600# a_3383_n655# a_3325_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X26 a_1261_n600# a_1061_n655# a_1003_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X27 a_n1835_n600# a_n2035_n655# a_n2093_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_XW23Q2 a_29_n964# a_n2351_n900# a_229_n900# a_n745_n964#
+ a_n1577_n900# a_2035_n900# a_803_n964# a_n2035_n964# a_n545_n900# a_1835_n964# a_1003_n900#
+ a_n229_n964# a_n1003_n964# a_287_n964# a_n2867_n900# a_2093_n964# a_487_n900# a_n29_n900#
+ a_2293_n900# a_1319_n964# a_n1835_n900# a_1061_n964# a_n2293_n964# a_n803_n900#
+ a_1519_n900# a_n2093_n900# a_n1519_n964# a_1261_n900# a_n487_n964# a_n1261_n964#
+ a_2609_n964# a_n1319_n900# a_545_n964# a_n287_n900# a_2351_n964# a_n1061_n900# a_1577_n964#
+ a_2809_n900# a_745_n900# a_n2809_n964# a_2551_n900# a_n2551_n964# w_n3067_n1197#
+ a_1777_n900# a_n2609_n900# a_n1777_n964#
X0 a_n2609_n900# a_n2809_n964# a_n2867_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1 a_1261_n900# a_1061_n964# a_1003_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X2 a_n1835_n900# a_n2035_n964# a_n2093_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X3 a_2809_n900# a_2609_n964# a_2551_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X4 a_n2351_n900# a_n2551_n964# a_n2609_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 a_n2093_n900# a_n2293_n964# a_n2351_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 a_n29_n900# a_n229_n964# a_n287_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X7 a_229_n900# a_29_n964# a_n29_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 a_n1319_n900# a_n1519_n964# a_n1577_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X9 a_2551_n900# a_2351_n964# a_2293_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 a_n545_n900# a_n745_n964# a_n803_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X11 a_n287_n900# a_n487_n964# a_n545_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 a_2293_n900# a_2093_n964# a_2035_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X13 a_n803_n900# a_n1003_n964# a_n1061_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X14 a_n1577_n900# a_n1777_n964# a_n1835_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X15 a_1519_n900# a_1319_n964# a_1261_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X16 a_n1061_n900# a_n1261_n964# a_n1319_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 a_1003_n900# a_803_n964# a_745_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X18 a_745_n900# a_545_n964# a_487_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X19 a_487_n900# a_287_n964# a_229_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X20 a_1777_n900# a_1577_n964# a_1519_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X21 a_2035_n900# a_1835_n964# a_1777_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HG2LSW a_n100_n205# a_100_n150# a_n292_n372#
+ a_n158_n150#
X0 a_100_n150# a_n100_n205# a_n158_n150# a_n292_n372# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N64HU4 a_3235_n255# a_n1861_n200# a_n1803_n255#
+ a_n3827_n422# a_n2777_n200# a_n1345_n255# a_n2719_n255# a_3635_n200# a_2261_n200#
+ a_n1403_n200# a_3177_n200# a_n2319_n200# a_1861_n255# a_2777_n255# a_1403_n255#
+ a_n887_n255# a_n945_n200# a_945_n255# a_2319_n255# a_n487_n200# a_n429_n255# a_1803_n200#
+ a_487_n255# a_2719_n200# a_1345_n200# a_n29_n200# a_n3693_n200# a_n2261_n255# a_n3635_n255#
+ a_887_n200# a_29_n255# a_n3177_n255# a_n3235_n200# a_429_n200#
X0 a_1345_n200# a_945_n255# a_887_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X1 a_n2319_n200# a_n2719_n255# a_n2777_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X2 a_n2777_n200# a_n3177_n255# a_n3235_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X3 a_2261_n200# a_1861_n255# a_1803_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X4 a_n945_n200# a_n1345_n255# a_n1403_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X5 a_3635_n200# a_3235_n255# a_3177_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X6 a_429_n200# a_29_n255# a_n29_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X7 a_1803_n200# a_1403_n255# a_1345_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X8 a_887_n200# a_487_n255# a_429_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X9 a_3177_n200# a_2777_n255# a_2719_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X10 a_n3235_n200# a_n3635_n255# a_n3693_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X11 a_n487_n200# a_n887_n255# a_n945_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X12 a_n1403_n200# a_n1803_n255# a_n1861_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X13 a_2719_n200# a_2319_n255# a_2261_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X14 a_n1861_n200# a_n2261_n255# a_n2319_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X15 a_n29_n200# a_n429_n255# a_n487_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RMXH5H a_803_n255# a_1261_n200# a_n1319_n200#
+ a_n287_n200# a_n229_n255# a_n1061_n200# a_287_n255# a_n1003_n255# a_745_n200# a_1319_n255#
+ a_n1711_n422# a_1061_n255# a_229_n200# a_n1577_n200# a_n1519_n255# a_n487_n255#
+ a_n545_n200# a_n1261_n255# a_545_n255# a_1003_n200# a_487_n200# a_n29_n200# a_29_n255#
+ a_n745_n255# a_n803_n200# a_1519_n200#
X0 a_487_n200# a_287_n255# a_229_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1261_n200# a_1061_n255# a_1003_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n29_n200# a_n229_n255# a_n287_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_229_n200# a_29_n255# a_n29_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X5 a_n545_n200# a_n745_n255# a_n803_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n287_n200# a_n487_n255# a_n545_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_1519_n200# a_1319_n255# a_1261_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X9 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_745_n200# a_545_n255# a_487_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_1003_n200# a_803_n255# a_745_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__res_high_po_0p69_XTGLEU a_282_n556# a_282_124# a_516_n556# a_48_124#
+ a_n186_124# a_n420_n556# a_n654_n556# a_516_124# a_48_n556# a_n784_n686# a_n420_124#
+ a_n654_124# a_n186_n556#
X0 a_n420_124# a_n420_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X1 a_48_124# a_48_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X2 a_282_124# a_282_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X3 a_516_124# a_516_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X4 a_n186_124# a_n186_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X5 a_n654_124# a_n654_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_TT9EEV a_n932_n420# a_1648_n420# a_n1648_n484#
+ a_1390_n420# a_n1390_n484# a_n616_n484# a_n1448_n420# a_674_n484# a_n1190_n420#
+ w_n1906_n717# a_n416_n420# a_874_n420# a_158_n484# a_358_n420# a_n874_n484# a_n1706_n420#
+ a_932_n484# a_100_n420# a_n674_n420# a_1132_n420# a_n358_n484# a_n1132_n484# a_416_n484#
+ a_n158_n420# a_n100_n484# a_616_n420# a_1448_n484# a_1190_n484#
X0 a_n416_n420# a_n616_n484# a_n674_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X1 a_n158_n420# a_n358_n484# a_n416_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X2 a_n1448_n420# a_n1648_n484# a_n1706_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=1.218 ps=8.98 w=4.2 l=1
X3 a_n1190_n420# a_n1390_n484# a_n1448_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X4 a_n674_n420# a_n874_n484# a_n932_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X5 a_n932_n420# a_n1132_n484# a_n1190_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X6 a_358_n420# a_158_n484# a_100_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X7 a_616_n420# a_416_n484# a_358_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X8 a_1648_n420# a_1448_n484# a_1390_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=1.218 pd=8.98 as=0.609 ps=4.49 w=4.2 l=1
X9 a_1132_n420# a_932_n484# a_874_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X10 a_874_n420# a_674_n484# a_616_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X11 a_1390_n420# a_1190_n484# a_1132_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X12 a_100_n420# a_n100_n484# a_n158_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BH2H9S a_n229_n1664# a_1061_n1664# a_n1835_n1600#
+ a_n2351_n1600# a_n1261_n1664# a_n1061_n1600# a_1319_n1664# a_1261_n1600# a_287_n1664#
+ a_n2035_n1664# a_2035_n1600# a_n1319_n1600# a_n1519_n1664# a_1519_n1600# a_487_n1600#
+ a_545_n1664# a_29_n1664# a_n487_n1664# a_n287_n1600# w_n2551_n1897# a_745_n1600#
+ a_2093_n1664# a_1577_n1664# a_803_n1664# a_n745_n1664# a_n1003_n1664# a_1003_n1600#
+ a_n545_n1600# a_n2293_n1664# a_n2093_n1600# a_n1777_n1664# a_2293_n1600# a_n1577_n1600#
+ a_1777_n1600# a_n29_n1600# a_1835_n1664# a_229_n1600# a_n803_n1600#
X0 a_n287_n1600# a_n487_n1664# a_n545_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X1 a_n1577_n1600# a_n1777_n1664# a_n1835_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X2 a_n29_n1600# a_n229_n1664# a_n287_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X3 a_2035_n1600# a_1835_n1664# a_1777_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X4 a_n1319_n1600# a_n1519_n1664# a_n1577_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X5 a_n2093_n1600# a_n2293_n1664# a_n2351_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=1
X6 a_745_n1600# a_545_n1664# a_487_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X7 a_n1835_n1600# a_n2035_n1664# a_n2093_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X8 a_1261_n1600# a_1061_n1664# a_1003_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X9 a_n545_n1600# a_n745_n1664# a_n803_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X10 a_229_n1600# a_29_n1664# a_n29_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X11 a_1003_n1600# a_803_n1664# a_745_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X12 a_n1061_n1600# a_n1261_n1664# a_n1319_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X13 a_n803_n1600# a_n1003_n1664# a_n1061_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X14 a_1777_n1600# a_1577_n1664# a_1519_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X15 a_1519_n1600# a_1319_n1664# a_1261_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X16 a_487_n1600# a_287_n1664# a_229_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X17 a_2293_n1600# a_2093_n1664# a_2035_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U a_n1861_n200# a_n1803_n255# a_n3369_n422#
+ a_n2777_n200# a_n1345_n255# a_n2719_n255# a_2261_n200# a_n1403_n200# a_3177_n200#
+ a_n2319_n200# a_1861_n255# a_2777_n255# a_1403_n255# a_n887_n255# a_n945_n200# a_945_n255#
+ a_2319_n255# a_n487_n200# a_n429_n255# a_1803_n200# a_487_n255# a_2719_n200# a_1345_n200#
+ a_n29_n200# a_n2261_n255# a_887_n200# a_29_n255# a_n3177_n255# a_n3235_n200# a_429_n200#
X0 a_1345_n200# a_945_n255# a_887_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X1 a_n2319_n200# a_n2719_n255# a_n2777_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X2 a_n2777_n200# a_n3177_n255# a_n3235_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X3 a_2261_n200# a_1861_n255# a_1803_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X4 a_n945_n200# a_n1345_n255# a_n1403_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X5 a_429_n200# a_29_n255# a_n29_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X6 a_1803_n200# a_1403_n255# a_1345_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X7 a_887_n200# a_487_n255# a_429_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X8 a_3177_n200# a_2777_n255# a_2719_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X9 a_n487_n200# a_n887_n255# a_n945_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X10 a_n1403_n200# a_n1803_n255# a_n1861_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X11 a_2719_n200# a_2319_n255# a_2261_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X12 a_n1861_n200# a_n2261_n255# a_n2319_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X13 a_n29_n200# a_n429_n255# a_n487_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
.ends

.subckt sky130_td_ip__opamp_hp avdd vout ibias vinn vinp dvdd ena dvss avss
Xsky130_fd_pr__pfet_g5v0d10v5_W75H7K_0 net4 avdd net5 net5 avdd net4 avdd net5 net5
+ net5 net5 net3 net5 net5 net3 net4 avdd avdd net5 net5 avdd net4 net3 avdd net5
+ net5 net5 avdd net3 net4 net5 avdd avdd net5 net5 avdd net3 net5 avdd net5 net5
+ net4 net5 net5 avdd net5 net3 avdd net5 net4 avdd net5 net5 avdd net4 net5 net5
+ net5 net4 net5 avdd net3 avdd net5 net3 net5 net4 avdd net3 avdd avdd net5 net5
+ net5 avdd net5 net5 avdd sky130_fd_pr__pfet_g5v0d10v5_W75H7K
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_15 avdd avdd m1_n3750_n668# net21 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_16 net5 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_WKXP7K_0 net3 m1_n592_3104# avdd vb2 vb2 net4 m1_n592_3104#
+ vb2 vb2 vb2 vb2 net3 vb2 vb2 net4 net4 net5 net5 vb2 vb2 m1_n592_3104# net3 net3
+ net5 vb2 vb2 vb2 m1_n592_3104# avdd net3 vb2 m1_n592_3104# net5 vb2 vb2 m1_n592_3104#
+ net3 avdd m1_n592_3104# vb2 vb2 net4 vb2 vb2 net5 vb2 avdd avdd avdd net4 net5 vb2
+ net4 net5 vb2 vb2 m1_n592_3104# net3 vb2 vb2 vb2 net3 vb2 m1_n592_3104# net3 m1_n592_3104#
+ vb2 net4 vb2 net4 net5 net4 net5 vb2 vb2 avdd vb2 net5 vb2 avdd vb2 vb2 sky130_fd_pr__pfet_g5v0d10v5_WKXP7K
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_17 m1_n3750_n668# avdd net35 avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_01v8_6H2JYD_0 dvss m1_n6583_10102# m1_n5758_10095# dvss sky130_fd_pr__nfet_01v8_6H2JYD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_0 ibias avss net33 m1_n3750_n668# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_HQ4STX_0 avdd vb2 vb2 avdd sky130_fd_pr__pfet_g5v0d10v5_HQ4STX
Xsky130_fd_pr__nfet_01v8_6H2JYD_1 dvss ena m1_n6583_10102# dvss sky130_fd_pr__nfet_01v8_6H2JYD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_1 net34 avss net31 m1_n3750_n668# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_2 m1_n3750_n668# avss avss net35 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_UKVZ7J_0 net29 avss net12 m1_n4692_n1074# avss m1_n4692_n1074#
+ m1_n4692_n1074# m1_n4692_n1074# avss avss net12 m1_n4692_n1074# m1_n4692_n1074#
+ avss m1_n4692_n1074# m1_n4692_n1074# avss avss net12 avss m1_n4692_n1074# net12
+ avss net12 m1_n4692_n1074# m1_n4692_n1074# avss m1_n4692_n1074# m1_n4692_n1074#
+ avss net29 avss net12 m1_n4692_n1074# net28 m1_n4692_n1074# m1_n4692_n1074# avss
+ net12 m1_n4692_n1074# avss m1_n4692_n1074# avss m1_n4692_n1074# m1_n4692_n1074#
+ net12 m1_n4692_n1074# net28 m1_n4692_n1074# avss avss net12 m1_n4692_n1074# m1_n4692_n1074#
+ sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_3 net6 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_USXRNR_0 avss net10 avss avss avss net6 net5 net10 net10
+ net10 net8 net5 avss net8 net10 net6 avss net10 m1_n592_3104# net6 net10 net6 net5
+ net10 m1_n592_3104# avss net10 avss sky130_fd_pr__nfet_g5v0d10v5_USXRNR
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_0 avdd avdd m1_n3750_n668# net3 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_4 net10 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_1 net18 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_5 vb3 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_2 avdd avdd m1_n3750_n668# vb1 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_6 m1_n4692_n1074# avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_AUMBFF_0 m1_n592_3104# m1_n592_3104# avdd vout avdd
+ vout avdd m1_n592_3104# m1_n592_3104# m1_n592_3104# vout m1_n592_3104# m1_n592_3104#
+ m1_n592_3104# m1_n592_3104# vout m1_n592_3104# m1_n592_3104# m1_n592_3104# avdd
+ avdd avdd avdd m1_n592_3104# m1_n592_3104# avdd vout avdd vout m1_n592_3104# m1_n592_3104#
+ vout avdd m1_n592_3104# vout avdd avdd avdd m1_n592_3104# avdd avdd m1_n592_3104#
+ vout vout m1_n592_3104# m1_n592_3104# vout avdd m1_n592_3104# m1_n592_3104# avdd
+ m1_n592_3104# m1_n592_3104# vout m1_n592_3104# avdd vout avdd m1_n592_3104# m1_n592_3104#
+ vout avdd m1_n592_3104# avdd m1_n592_3104# m1_n592_3104# m1_n592_3104# vout avdd
+ vout sky130_fd_pr__pfet_g5v0d10v5_AUMBFF
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_3 vb5 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_7 net33 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__diode_pw2nd_05v5_25PWK4_0 dvss ena sky130_fd_pr__diode_pw2nd_05v5_25PWK4
Xsky130_fd_pr__pfet_g5v0d10v5_QL2RRT_0 vinn vinn net1 vinp net1 vtailp vinp vtailp
+ vinp vinn vtailp avdd vinn vtailp vinn avdd vinn vinp net2 avdd vinn avdd vtailp
+ vtailp vinp net1 vtailp vinn net1 vinp net2 vtailp vtailp vinp net2 vinn vinp vinp
+ vinp net2 net1 vtailp vinn net2 vinn net2 avdd vinp vtailp vinn vtailp net1 vtailp
+ vinp sky130_fd_pr__pfet_g5v0d10v5_QL2RRT
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_4 net13 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_8 net20 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QL2RRT_1 vinp vinp net2 vinn net2 vtailp vinn vtailp
+ vinn vinp vtailp avdd vinp vtailp vinp avdd vinp vinn net1 avdd vinp avdd vtailp
+ vtailp vinn net2 vtailp vinp net2 vinn net1 vtailp vtailp vinn net1 vinp vinn vinn
+ vinn net1 net2 vtailp vinp net1 vinp net1 avdd vinn vtailp vinp vtailp net2 vtailp
+ vinn sky130_fd_pr__pfet_g5v0d10v5_QL2RRT
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_5 avdd avdd m1_n3667_4379# enab_avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_9 net31 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_7 avdd avdd m1_n3750_n668# m1_791_7588# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_6 avdd avdd m1_n3750_n668# vb2 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_01v8_U4BBJH_1 m1_n6583_10102# dvdd ena dvdd sky130_fd_pr__pfet_01v8_U4BBJH
Xsky130_fd_pr__pfet_01v8_U4BBJH_0 m1_n5758_10095# dvdd m1_n6583_10102# dvdd sky130_fd_pr__pfet_01v8_U4BBJH
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_8 m1_180_4838# avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_9 net4 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_QTY6KC_0 m1_18668_3467# m1_180_4838# m1_18668_3467#
+ avdd avdd avdd m1_18668_3467# avdd m1_18668_3467# avdd avdd m1_180_4838# m1_180_4838#
+ m1_18668_3467# m1_18668_3467# m1_18668_3467# m1_180_4838# avdd avdd m1_180_4838#
+ avdd avdd m1_18668_3467# m1_180_4838# m1_18668_3467# avdd sky130_fd_pr__pfet_g5v0d10v5_QTY6KC
Xsky130_fd_pr__nfet_g5v0d10v5_B3XH3Z_0 vtailn avss vb1 avss net12 vb3 vb3 vb3 net29
+ avss vtailn avss net12 vb1 vb3 avss net12 vb3 vb3 net12 net28 avss vtailn vb3 vb3
+ vtailn net12 m1_n4692_n1074# vb3 avss avss vb3 vb3 net12 vb1 vb3 vtailn avss vb3
+ vtailn avss vb3 avss vtailn m1_n4692_n1074# vb3 vb3 net28 vb3 net12 vb3 vb3 vtailn
+ vb3 vtailn vb3 vb3 net12 net29 m1_n4692_n1074# vb3 vb3 sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_10 net12 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QTY6H6_0 avdd net22 net22 avdd net22 avdd m1_n3445_8429#
+ avdd net22 avdd net22 avdd net22 m1_n3445_8429# m1_n3445_8429# net22 net22 net22
+ m1_n3445_8429# net32 avdd net22 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5_QTY6H6
Xsky130_fd_pr__nfet_g5v0d10v5_U73S5M_0 vout vout net8 net8 net8 avss avss vout avss
+ net8 net8 avss vout vout avss net8 net8 net8 net8 net8 net8 avss avss net8 vout
+ avss net8 vout vout avss net8 net8 avss net8 avss avss vout vout net8 avss net8
+ net8 vout net8 net8 net8 net8 net8 net8 net8 avss vout net8 avss avss net8 net8
+ net8 avss vout vout net8 avss net8 vout avss avss vout avss avss sky130_fd_pr__nfet_g5v0d10v5_U73S5M
Xsky130_fd_pr__pfet_g5v0d10v5_PP2RNK_0 vb2 vb1 vtailp avdd vb2 avdd m1_791_7588# vb2
+ vb2 m1_791_7588# avdd vb2 m1_791_7588# vb2 vb2 vb2 vb1 vb2 m1_791_7588# m1_791_7588#
+ vtailp avdd vb2 vb1 vb2 vb2 vtailp m1_791_7588# m1_3549_9621# avdd vtailp vb2 vb2
+ vb2 vtailp vb2 vtailp vb2 m1_791_7588# vb2 vtailp vtailp vb2 m1_791_7588# vb2 avdd
+ vtailp m1_3549_9621# avdd avdd sky130_fd_pr__pfet_g5v0d10v5_PP2RNK
Xsky130_fd_pr__nfet_g5v0d10v5_79TVLH_0 vtailn net4 vtailn vinn vinp net4 net4 vtailn
+ vinn vtailn vinp vtailn vinn vinn vinn avss vinp vtailn vinp net3 vinn avss vinp
+ vtailn vtailn vinn vinp vinp net4 net4 vtailn vinn vinn vtailn net3 vtailn vinn
+ vinp net3 net3 avss vinp net4 vinp vtailn vinp vinn net3 net3 vinp avss avss vtailn
+ vinn sky130_fd_pr__nfet_g5v0d10v5_79TVLH
Xsky130_fd_pr__nfet_g5v0d10v5_2B7385_0 avss avss m1_n5910_1250# avss m1_n5910_1250#
+ m1_n5910_1250# m1_n5910_1250# m1_n5910_1250# avss avss m1_n5910_1250# avss avss
+ avss m1_n5910_1250# avss vtailn vtailn m1_n5910_1250# m1_n5910_1250# m1_n5910_1250#
+ vtailn m1_n5910_1250# m1_n5910_1250# m1_n5910_1250# avss vtailn vtailn avss m1_n5910_1250#
+ m1_n5910_1250# avss m1_n5910_1250# avss vtailn vtailn m1_n5910_1250# m1_n5910_1250#
+ sky130_fd_pr__nfet_g5v0d10v5_2B7385
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_11 net2 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_79TVLH_1 vtailn net3 vtailn vinp vinn net3 net3 vtailn
+ vinp vtailn vinn vtailn vinp vinp vinp avss vinn vtailn vinn net4 vinp avss vinn
+ vtailn vtailn vinp vinn vinn net3 net3 vtailn vinp vinp vtailn net4 vtailn vinp
+ vinn net4 net4 avss vinn net3 vinn vtailn vinn vinp net4 net4 vinn avss avss vtailn
+ vinp sky130_fd_pr__nfet_g5v0d10v5_79TVLH
Xsky130_fd_pr__nfet_g5v0d10v5_NT3TPY_0 m1_n5758_10095# net35 avss avss avss avss net35
+ avss avss m1_n3667_4379# m1_n6583_10102# avss m1_n6583_10102# m1_n5758_10095# sky130_fd_pr__nfet_g5v0d10v5_NT3TPY
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_12 net1 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_5X2ZTR_0 vb2 vb7 vb7 vb7 avss net16 avss vb6 net24 vb7
+ avss vb7 avss net16 vb7 vb6 avss vb7 avss net25 net16 net24 avss vb7 vb6 vb6 vb7
+ vb7 net25 net16 vb2 vb7 vb7 avss net24 net16 vb7 vb2 vb8 vb7 vb7 avss net25 avss
+ vb7 m1_180_4838# net24 avss avss net25 vb7 vb7 vb7 vb2 vb7 m1_180_4838# avss avss
+ vb7 vb7 net25 net24 vb7 vb7 vb7 m1_180_4838# m1_180_4838# vb7 net25 vb7 vb7 vb7
+ net24 vb2 vb7 vb7 vb7 vb7 net16 vb7 vb6 m1_180_4838# sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR
Xsky130_fd_pr__nfet_g5v0d10v5_WK95DB_0 avss net18 vb3 vb3 vb3 vtailn vtailn vb3 vb3
+ net18 net18 vb3 vb3 vtailn vb3 avss net18 avss avss avss net18 vtailn sky130_fd_pr__nfet_g5v0d10v5_WK95DB
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_13 vb7 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14 vinp avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_15 m1_n5910_1250# avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_3QL9S5_0 enab_avdd m1_12266_11884# avdd net21 sky130_fd_pr__pfet_g5v0d10v5_3QL9S5
Xsky130_fd_pr__nfet_g5v0d10v5_PGZBW9_0 net6 net6 net1 net1 avss net6 avss net6 net6
+ avss net6 net6 net6 avss avss net6 net2 net6 avss net6 avss avss net6 net6 net1
+ avss net6 net1 net6 net6 net2 avss avss net6 net6 net2 avss net2 net6 net1 avss
+ net6 net6 net6 net2 net6 net2 avss avss avss avss net1 avss net6 sky130_fd_pr__nfet_g5v0d10v5_PGZBW9
Xsky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD_1 avdd net35 avdd net35 avdd net35 avdd avdd
+ avdd net35 m1_n3667_4379# avdd avdd avdd m1_n3667_4379# m1_n3667_4379# m1_n3667_4379#
+ m1_n3667_4379# m1_n3667_4379# net35 avdd net35 sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_16 vb8 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_3QL9S5_1 enab_avdd net22 avdd net32 sky130_fd_pr__pfet_g5v0d10v5_3QL9S5
Xsky130_fd_pr__pfet_g5v0d10v5_QSKB8C_0 vb6 vb6 avdd vb3 vb6 vb5 vb6 m1_n4692_n1074#
+ m1_n4692_n1074# vb6 vb6 net13 m1_25484_9858# vb3 vb6 avdd vb6 net10 m1_25484_9858#
+ vb6 vb6 m1_n4692_n1074# vb6 vb6 net13 vb6 vb6 avdd m1_25484_9858# avdd avdd vb6
+ m1_25484_9858# m1_23420_9858# vb6 vb6 m1_n4692_n1074# vb6 vb6 avdd avdd vb6 avdd
+ m1_23420_9858# avdd net10 vb6 vb6 avdd vb6 net13 m1_n4692_n1074# avdd vb6 vb6 vb6
+ avdd m1_25484_9858# vb6 vb6 m1_25484_9858# m1_n4692_n1074# vb3 avdd net10 avdd vb6
+ vb5 vb6 vb5 m1_n4692_n1074# m1_23420_9858# vb6 vb6 vb6 net10 vb3 vb6 sky130_fd_pr__pfet_g5v0d10v5_QSKB8C
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_17 net16 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QRKB8C_0 vb5 vb5 avdd m1_23420_9858# vb5 avdd avdd vb5
+ vb5 avdd vb5 avdd avdd net13 vb5 vb5 avdd m1_25484_9858# avdd avdd avdd m1_25484_9858#
+ vb5 avdd avdd vb5 vb5 avdd vb5 vb5 m1_23420_9858# avdd avdd avdd m1_23420_9858#
+ m1_25484_9858# vb5 vb5 avdd vb5 avdd avdd vb5 net13 vb5 vb5 net13 avdd net13 vb5
+ vb5 vb5 vb5 avdd vb5 vb5 avdd m1_25484_9858# avdd vb5 m1_25484_9858# vb5 vb5 avdd
+ vb5 avdd vb5 avdd avdd vb5 vb5 m1_25484_9858# m1_23420_9858# vb5 sky130_fd_pr__pfet_g5v0d10v5_QRKB8C
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18 vinn avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__cap_mim_m3_1_Z5XS7R_1 net8 m1_n592_3104# m1_32750_1661# net8 m1_32495_1140#
+ m1_32495_1140# m1_n592_3104# net8 m1_32495_1140# m1_32750_1661# m1_32750_1661# m1_n592_3104#
+ sky130_fd_pr__cap_mim_m3_1_Z5XS7R
Xsky130_fd_pr__pfet_g5v0d10v5_EVM3FM_0 vb2 vb2 vb2 m1_n5910_1250# vb2 vb2 vtailp vb2
+ avdd vb2 vtailp vb2 avdd m1_n5910_1250# avdd avdd vtailp m1_n5910_1250# m1_n5910_1250#
+ avdd vtailp vtailp sky130_fd_pr__pfet_g5v0d10v5_EVM3FM
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_19 avss avss enab_avdd m1_n3667_4379# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_DL2ZHN_0 net16 vb8 vb8 vb8 avss vb8 net24 avss avss
+ vb8 vb8 avss vb8 net25 net16 vb8 vb8 avss avss avss vb8 vb8 net16 net24 vb8 vb8
+ avss avss net16 vb8 vb8 avss avss vb8 net25 net25 vb8 vb8 avss net16 vb8 net24 avss
+ vb8 avss avss vb8 vb8 net24 vb8 net16 vb8 net25 avss vb8 avss avss avss vb8 vb8
+ net24 vb8 avss avss vb8 vb8 avss avss net24 avss vb8 vb8 vb8 avss avss net25 net25
+ avss sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN
Xsky130_fd_pr__pfet_g5v0d10v5_Q46EE6_0 m1_n3445_8429# m1_12266_11884# m1_12266_11884#
+ avdd net21 m1_12266_11884# m1_n3445_8429# net32 avdd m1_n3445_8429# avdd avdd m1_12266_11884#
+ m1_n3445_8429# avdd net32 m1_12266_11884# vb7 vb7 m1_12266_11884# avdd m1_12266_11884#
+ vb7 vb7 m1_12266_11884# avdd m1_12266_11884# avdd vb7 m1_12266_11884# sky130_fd_pr__pfet_g5v0d10v5_Q46EE6
Xsky130_fd_pr__nfet_g5v0d10v5_UGZTXE_0 vb3 vb3 net6 net8 net1 avss vb3 net2 vb3 vb3
+ net1 vb3 vb3 vb3 avss net2 avss vb3 net6 vb3 net8 vb3 avss net2 vb3 vb3 net8 net1
+ avss net6 vb3 vb3 net6 net2 net1 vb3 vb3 avss net8 vb3 avss net6 vb3 net6 net1 avss
+ vb3 vb3 net8 vb3 net8 net6 vb3 net2 net2 net8 net1 vb3 sky130_fd_pr__nfet_g5v0d10v5_UGZTXE
Xsky130_fd_pr__pfet_g5v0d10v5_XW23Q2_0 vb1 m1_791_7588# m1_3549_9621# vb1 avdd avdd
+ vb1 vb1 avdd vb1 avdd vb1 vb1 vb1 avdd vb1 avdd avdd m1_791_7588# vb1 m1_791_7588#
+ vb1 vb1 m1_791_7588# avdd avdd vb1 m1_791_7588# vb1 vb1 avdd m1_791_7588# vb1 m1_3549_9621#
+ vb1 avdd vb1 avdd m1_791_7588# avdd avdd vb1 avdd m1_791_7588# avdd vb1 sky130_fd_pr__pfet_g5v0d10v5_XW23Q2
Xsky130_fd_pr__nfet_g5v0d10v5_HG2LSW_0 vb3 vb3 avss avss sky130_fd_pr__nfet_g5v0d10v5_HG2LSW
Xsky130_fd_pr__nfet_g5v0d10v5_N64HU4_0 avss avss avss avss ibias net33 net33 avss
+ net20 net20 net20 net34 net33 net33 net33 net33 net21 net33 net33 net20 net33 net21
+ net33 net21 net20 net21 avss avss avss net21 net33 net33 net34 net20 sky130_fd_pr__nfet_g5v0d10v5_N64HU4
Xsky130_fd_pr__nfet_g5v0d10v5_RMXH5H_0 m1_18790_1436# avss net10 net10 avss m1_18790_1436#
+ m1_18790_1436# net10 avss avss avss m1_18790_1436# avss avss avss net10 m1_18790_1436#
+ net10 m1_18790_1436# m1_18790_1436# m1_18790_1436# avss avss net10 net10 avss sky130_fd_pr__nfet_g5v0d10v5_RMXH5H
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_10 net32 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__res_high_po_0p69_XTGLEU_0 m1_32032_n77# m1_32750_1661# avss m1_32495_1140#
+ vout m1_32032_n77# avss avss m1_32268_124# avss vout avss m1_32268_124# sky130_fd_pr__res_high_po_0p69_XTGLEU
Xsky130_fd_pr__pfet_g5v0d10v5_TT9EEV_0 net5 avdd avdd net8 m1_180_4838# m1_180_4838#
+ net5 m1_180_4838# net6 avdd net5 net8 avdd avdd m1_180_4838# avdd m1_180_4838# net5
+ net6 m1_n592_3104# m1_180_4838# m1_180_4838# avdd net6 m1_180_4838# m1_n592_3104#
+ avdd m1_180_4838# sky130_fd_pr__pfet_g5v0d10v5_TT9EEV
Xsky130_fd_pr__pfet_g5v0d10v5_BH2H9S_0 net18 net18 vtailp avdd net18 avdd net18 vtailp
+ net18 net18 avdd vtailp net18 avdd avdd net18 net18 net18 net18 avdd vtailp avdd
+ net18 net18 net18 net18 avdd avdd avdd avdd net18 avdd avdd vtailp avdd net18 net18
+ vtailp sky130_fd_pr__pfet_g5v0d10v5_BH2H9S
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_11 net22 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_NMXZ6U_0 net20 net31 avss net20 net31 net31 avss avss
+ avss avss net31 avss net31 net31 net20 net31 net31 avss net31 net20 net31 net20
+ avss net34 net31 net20 net31 avss avss avss sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_12 avdd avdd m1_n3750_n668# vb6 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_14 avdd avdd m1_n3750_n668# m1_n3445_8429# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13 avdd avdd m1_n3750_n668# m1_n592_3104# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_HTFGEA a_n150_n150# a_n48_n48#
X0 a_n150_n150# a_n48_n48# sky130_fd_pr__diode_pw2nd_05v5 perim=1.92e+06 area=2.304e+11
.ends

.subckt sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X2 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X3 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6 w_n387_n462# a_29_n261# a_n129_n261# a_n29_n164#
+ a_n187_n164# a_129_n164#
X0 a_129_n164# a_29_n261# a_n29_n164# w_n387_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n164# a_n129_n261# a_n187_n164# w_n387_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HRGQF2 a_n321_n622# a_n29_n400# a_n187_n400#
+ a_129_n400# a_29_n488# a_n129_n488#
X0 a_n29_n400# a_n129_n488# a_n187_n400# a_n321_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_129_n400# a_29_n488# a_n29_n400# a_n321_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U62SY6 a_n187_n64# w_n387_n362# a_129_n64# a_29_n161#
+ a_n129_n161# a_n29_n64#
X0 a_129_n64# a_29_n161# a_n29_n64# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n64# a_n129_n161# a_n187_n64# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4 a_n242_n622# a_50_n400# a_n108_n400# a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n242_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6 a_n108_n164# a_n50_n261# w_n308_n462#
+ a_50_n164#
X0 a_50_n164# a_n50_n261# a_n108_n164# w_n308_n462# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ3N a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt isolated_switch on vss out in vdd
Xsky130_fd_pr__pfet_g5v0d10v5_U6V9Y6_0 vdd onb onb m1_1166_n2330# out out sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6
Xsky130_fd_pr__nfet_g5v0d10v5_HRGQF2_0 vss m1_1166_n2330# out out onp onp sky130_fd_pr__nfet_g5v0d10v5_HRGQF2
Xsky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 onb vdd onb on on vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM1 vss in m1_1166_n2330# m1_1166_n2330# onp onp sky130_fd_pr__nfet_g5v0d10v5_HRGQF2
XXM3 vss in in onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
XXM4 vdd onb onb in m1_1166_n2330# m1_1166_n2330# sky130_fd_pr__pfet_g5v0d10v5_U6V9Y6
XXM5 vss m1_1166_n2330# m1_1166_n2330# onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
XXM6 m1_1166_n2330# onp vdd m1_1166_n2330# sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
XXM7 onp vdd onp onb onb vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
Xsky130_fd_pr__nfet_g5v0d10v5_UNEQ3N_0 vss vss m1_1166_n2330# onb sky130_fd_pr__nfet_g5v0d10v5_UNEQ3N
XXM8 onp vss vss onb sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXD1 vss on sky130_fd_pr__diode_pw2nd_05v5_FT76RK
Xsky130_fd_pr__nfet_g5v0d10v5_MJGQJ4_0 vss m1_1166_n2330# m1_1166_n2330# onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
Xsky130_fd_pr__nfet_g5v0d10v5_MJGQJ4_1 vss out out onb sky130_fd_pr__nfet_g5v0d10v5_MJGQJ4
Xsky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_0 in onp vdd in sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
Xsky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_1 m1_1166_n2330# onp vdd m1_1166_n2330# sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
Xsky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6_2 out onp vdd out sky130_fd_pr__pfet_g5v0d10v5_U6Z9Y6
XXM10 onb vss vss on sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
.ends

.subckt analog_mux_sel1v8 selA dvdd out inA inB avdd avss dvss
Xsky130_fd_pr__diode_pw2nd_05v5_HTFGEA_0 dvss selA sky130_fd_pr__diode_pw2nd_05v5_HTFGEA
Xsky130_fd_sc_hvl__inv_2_0 isolated_switch_1/on dvss dvss avdd avdd isolated_switch_2/on
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 selA dvdd dvss dvss avdd avdd isolated_switch_1/on
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xisolated_switch_1 isolated_switch_1/on avss inA out avdd isolated_switch
Xisolated_switch_2 isolated_switch_2/on avss inB out avdd isolated_switch
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6 a_n29_n400# a_n187_n400# a_n345_n400#
+ a_29_n497# a_n129_n497# a_187_n497# a_129_n400# a_n503_n400# a_n287_n497# w_n861_n697#
+ a_287_n400# a_n661_n400# a_345_n497# a_n445_n497# a_445_n400# a_503_n497# a_n603_n497#
+ a_603_n400#
X0 a_n503_n400# a_n603_n497# a_n661_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_n29_n400# a_n129_n497# a_n187_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n497# a_445_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n187_n400# a_n287_n497# a_n345_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_287_n400# a_187_n497# a_129_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_n345_n400# a_n445_n497# a_n503_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X6 a_129_n400# a_29_n497# a_n29_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_445_n400# a_345_n497# a_287_n400# w_n861_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ a_n287_n488# a_345_n488# a_n29_n400# a_n187_n400#
+ a_n445_n488# a_503_n488# a_n345_n400# a_n603_n488# a_129_n400# a_n503_n400# a_287_n400#
+ a_n661_n400# a_445_n400# a_29_n488# a_n129_n488# a_603_n400# a_187_n488# a_n795_n622#
X0 a_n503_n400# a_n603_n488# a_n661_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_n29_n400# a_n129_n488# a_n187_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n488# a_445_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n187_n400# a_n287_n488# a_n345_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X4 a_287_n400# a_187_n488# a_129_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_n345_n400# a_n445_n488# a_n503_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X6 a_129_n400# a_29_n488# a_n29_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_445_n400# a_345_n488# a_287_n400# a_n795_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__diode_pd2nw_11v0_K4SERG a_n45_n45# w_n243_n243#
X0 a_n45_n45# w_n243_n243# sky130_fd_pr__diode_pd2nw_11v0 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6 a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt level_shifter_ad AVDD LO_B LO HI HI_B AVSS
XXM25 HI AVDD AVDD HI_B sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM1 HI_B HI AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM2 HI AVSS AVSS LO_B sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM21 AVSS AVSS HI_B LO sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
.ends

.subckt sky130_fd_pr__diode_pw2nd_11v0_FT76RJ a_n181_n181# a_n45_n45#
X0 a_n181_n181# a_n45_n45# sky130_fd_pr__diode_pw2nd_11v0 perim=1.8e+06 area=2.025e+11
.ends

.subckt power_gating_ad ENA STDBY IBIAS EG_AVDD EG_AVSS SG_AVDD SG_AVSS EG_IBIAS XIN
+ ENA_B STDBY_B AVSS AVDD
XXM25 AVDD EG_AVDD AVDD level_shifter_ad_0/HI_B level_shifter_ad_0/HI_B level_shifter_ad_0/HI_B
+ EG_AVDD EG_AVDD level_shifter_ad_0/HI_B AVDD AVDD AVDD level_shifter_ad_0/HI_B level_shifter_ad_0/HI_B
+ EG_AVDD level_shifter_ad_0/HI_B level_shifter_ad_0/HI_B AVDD sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6
XXM1 AVDD SG_AVDD AVDD level_shifter_ad_1/HI level_shifter_ad_1/HI level_shifter_ad_1/HI
+ SG_AVDD SG_AVDD level_shifter_ad_1/HI AVDD AVDD AVDD level_shifter_ad_1/HI level_shifter_ad_1/HI
+ SG_AVDD level_shifter_ad_1/HI level_shifter_ad_1/HI AVDD sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6
Xsky130_fd_pr__nfet_g5v0d10v5_CPEQJZ_0 level_shifter_ad_0/HI level_shifter_ad_0/HI
+ EG_AVSS AVSS level_shifter_ad_0/HI level_shifter_ad_0/HI EG_AVSS level_shifter_ad_0/HI
+ AVSS AVSS EG_AVSS EG_AVSS AVSS level_shifter_ad_0/HI level_shifter_ad_0/HI EG_AVSS
+ level_shifter_ad_0/HI AVSS sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ
Xsky130_fd_pr__nfet_g5v0d10v5_CPEQJZ_1 level_shifter_ad_1/HI_B level_shifter_ad_1/HI_B
+ SG_AVSS AVSS level_shifter_ad_1/HI_B level_shifter_ad_1/HI_B SG_AVSS level_shifter_ad_1/HI_B
+ AVSS AVSS SG_AVSS SG_AVSS AVSS level_shifter_ad_1/HI_B level_shifter_ad_1/HI_B SG_AVSS
+ level_shifter_ad_1/HI_B AVSS sky130_fd_pr__nfet_g5v0d10v5_CPEQJZ
Xsky130_fd_pr__diode_pd2nw_11v0_K4SERG_0 XIN AVDD sky130_fd_pr__diode_pd2nw_11v0_K4SERG
Xlevel_shifter_ad_0 AVDD ENA_B ENA level_shifter_ad_0/HI level_shifter_ad_0/HI_B AVSS
+ level_shifter_ad
Xlevel_shifter_ad_1 AVDD STDBY_B STDBY level_shifter_ad_1/HI level_shifter_ad_1/HI_B
+ AVSS level_shifter_ad
Xsky130_fd_pr__diode_pw2nd_11v0_FT76RJ_0 AVSS XIN sky130_fd_pr__diode_pw2nd_11v0_FT76RJ
Xsky130_fd_pr__pfet_g5v0d10v5_KL7ZY6_0 IBIAS EG_IBIAS IBIAS level_shifter_ad_0/HI_B
+ level_shifter_ad_0/HI_B level_shifter_ad_0/HI_B EG_IBIAS EG_IBIAS level_shifter_ad_0/HI_B
+ AVDD IBIAS IBIAS level_shifter_ad_0/HI_B level_shifter_ad_0/HI_B EG_IBIAS level_shifter_ad_0/HI_B
+ level_shifter_ad_0/HI_B IBIAS sky130_fd_pr__pfet_g5v0d10v5_KL7ZY6
.ends

.subckt sky130_fd_pr__nfet_01v8_HNLS5R a_n273_422# a_n413_n400# a_255_n400# a_351_n400#
+ a_n129_n400# a_63_n400# a_n225_n400# a_n321_n400# a_111_422# a_207_n488# a_n33_n400#
+ a_n369_n488# a_303_422# a_15_n488# a_n81_422# a_n177_n488# a_159_n400# a_n515_n574#
X0 a_n225_n400# a_n273_422# a_n321_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1 a_63_n400# a_15_n488# a_n33_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2 a_n129_n400# a_n177_n488# a_n225_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3 a_n33_n400# a_n81_422# a_n129_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X4 a_351_n400# a_303_422# a_255_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X5 a_255_n400# a_207_n488# a_159_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X6 a_n321_n400# a_n369_n488# a_n413_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X7 a_159_n400# a_111_422# a_63_n400# a_n515_n574# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt level_shifter_dd DVDD LO LO_B DVSS
XXM27 DVDD LO_B DVDD LO sky130_fd_pr__pfet_01v8_XGS3BL
XXM18 DVSS LO LO_B DVSS sky130_fd_pr__nfet_01v8_648S5X
.ends

.subckt sky130_fd_pr__pfet_01v8_XGNZDL a_n413_n400# a_111_431# a_255_n400# a_207_n497#
+ a_351_n400# a_n369_n497# a_303_431# a_n129_n400# a_63_n400# a_n225_n400# a_15_n497#
+ a_n81_431# a_n177_n497# a_n273_431# a_n321_n400# w_n551_n619# a_n33_n400# a_159_n400#
X0 a_n129_n400# a_n177_n497# a_n225_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1 a_n33_n400# a_n81_431# a_n129_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2 a_351_n400# a_303_431# a_255_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3 a_255_n400# a_207_n497# a_159_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X4 a_n321_n400# a_n369_n497# a_n413_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X5 a_159_n400# a_111_431# a_63_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X6 a_n225_n400# a_n273_431# a_n321_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X7 a_63_n400# a_15_n497# a_n33_n400# w_n551_n619# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
.ends

.subckt power_gating_dd ENA ENA_B STDBY STDBY_B SG_DVSS SG_DVDD DOUT DVDD DVSS
XXM18 STDBY_B SG_DVSS DVSS SG_DVSS DVSS DVSS SG_DVSS DVSS STDBY_B STDBY_B SG_DVSS
+ STDBY_B STDBY_B STDBY_B STDBY_B STDBY_B SG_DVSS DVSS sky130_fd_pr__nfet_01v8_HNLS5R
Xsky130_fd_pr__nfet_01v8_HNLS5R_0 STDBY DOUT DVSS DOUT DVSS DVSS DOUT DVSS STDBY STDBY
+ DOUT STDBY STDBY STDBY STDBY STDBY DOUT DVSS sky130_fd_pr__nfet_01v8_HNLS5R
Xlevel_shifter_dd_0 DVDD ENA ENA_B DVSS level_shifter_dd
Xlevel_shifter_dd_1 DVDD STDBY STDBY_B DVSS level_shifter_dd
Xsky130_fd_pr__pfet_01v8_XGNZDL_0 DVDD STDBY SG_DVDD STDBY DVDD STDBY STDBY SG_DVDD
+ SG_DVDD DVDD STDBY STDBY STDBY STDBY SG_DVDD DVDD DVDD DVDD sky130_fd_pr__pfet_01v8_XGNZDL
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MPZGNS m3_n1686_n9840# c1_n1646_n9800#
X0 c1_n1646_n9800# m3_n1686_n9840# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X1 c1_n1646_n9800# m3_n1686_n9840# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X2 c1_n1646_n9800# m3_n1686_n9840# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X3 c1_n1646_n9800# m3_n1686_n9840# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X4 c1_n1646_n9800# m3_n1686_n9840# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X5 c1_n1646_n9800# m3_n1686_n9840# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
.ends

.subckt power_gating DOUT SG_AVDD EG_IBIAS SG_DVDD AVDD EG_AVDD ENA SG_DVSS SG_AVSS
+ STDBY EG_AVSS XIN li_4587_n15047# AVSS DVDD IBIAS DVSS
Xpower_gating_ad_1 ENA STDBY IBIAS EG_AVDD EG_AVSS SG_AVDD SG_AVSS EG_IBIAS XIN power_gating_dd_0/ENA_B
+ power_gating_dd_0/STDBY_B AVSS AVDD power_gating_ad
Xpower_gating_dd_0 ENA power_gating_dd_0/ENA_B STDBY power_gating_dd_0/STDBY_B SG_DVSS
+ SG_DVDD DOUT DVDD DVSS power_gating_dd
XXC3 AVSS AVDD sky130_fd_pr__cap_mim_m3_1_MPZGNS
XXC4 DVSS DVDD sky130_fd_pr__cap_mim_m3_1_MPZGNS
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_33YP5M a_214_n832# a_214_400# a_n284_400#
+ a_48_n832# a_n118_400# a_n284_n832# a_n414_n962# a_n118_n832# a_48_400#
X0 a_214_400# a_214_n832# a_n414_n962# sky130_fd_pr__res_xhigh_po_0p35 l=4.16
X1 a_n284_400# a_n284_n832# a_n414_n962# sky130_fd_pr__res_xhigh_po_0p35 l=4.16
X2 a_48_400# a_48_n832# a_n414_n962# sky130_fd_pr__res_xhigh_po_0p35 l=4.16
X3 a_n118_400# a_n118_n832# a_n414_n962# sky130_fd_pr__res_xhigh_po_0p35 l=4.16
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_METDPQ a_546_n2036# a_n284_1604# a_n118_1604#
+ a_n284_n2036# a_n616_n2036# a_380_1604# a_n118_n2036# a_n616_1604# a_214_1604# a_380_n2036#
+ a_n746_n2166# a_48_1604# a_n450_n2036# a_214_n2036# a_546_1604# a_48_n2036# a_n450_1604#
X0 a_n118_1604# a_n118_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X1 a_n616_1604# a_n616_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X2 a_380_1604# a_380_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X3 a_546_1604# a_546_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X4 a_n450_1604# a_n450_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X5 a_n284_1604# a_n284_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X6 a_48_1604# a_48_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
X7 a_214_1604# a_214_n2036# a_n746_n2166# sky130_fd_pr__res_xhigh_po_0p35 l=16.2
.ends

.subckt sky130_fd_pr__pfet_01v8_6QYSWZ a_n88_n100# w_n226_n319# a_30_n100# a_n33_n197#
X0 a_30_n100# a_n33_n197# a_n88_n100# w_n226_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_723X3M a_20_n100# a_n78_n100# a_n33_n188# a_n180_n274#
X0 a_20_n100# a_n33_n188# a_n78_n100# a_n180_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.2
.ends

.subckt schmitt_trigger_pullmid SG_DVDD AIN DOUT SG_DVSS
Xsky130_fd_pr__res_xhigh_po_0p35_33YP5M_0 SG_DVDD m1_4000_3180# m1_3670_3180# m1_3830_1980#
+ m1_3670_3180# m1_3280_n190# SG_DVSS m1_3830_1980# m1_4000_3180# sky130_fd_pr__res_xhigh_po_0p35_33YP5M
XXR2 m1_4000_n1770# SG_DVSS m1_3280_n190# m1_4000_n1770# m1_3830_n540# m1_3670_n1770#
+ SG_DVSS m1_3670_n1770# m1_3830_n540# sky130_fd_pr__res_xhigh_po_0p35_33YP5M
XXR3 m1_3110_n1770# m1_2280_1870# m1_2620_1870# m1_2450_n1770# m1_2120_n1770# m1_2950_1870#
+ m1_2450_n1770# AIN m1_2950_1870# m1_3110_n1770# SG_DVSS m1_2620_1870# m1_2120_n1770#
+ m1_2780_n1770# m1_3280_n190# m1_2780_n1770# m1_2280_1870# sky130_fd_pr__res_xhigh_po_0p35_METDPQ
XXM3 m1_3799_1180# SG_DVDD DOUT AIN sky130_fd_pr__pfet_01v8_6QYSWZ
XXM4 m1_3800_300# DOUT AIN SG_DVSS sky130_fd_pr__nfet_01v8_723X3M
XXM5 SG_DVDD SG_DVDD m1_3799_1180# AIN sky130_fd_pr__pfet_01v8_6QYSWZ
XXM6 SG_DVSS m1_3800_300# AIN SG_DVSS sky130_fd_pr__nfet_01v8_723X3M
XXM7 m1_3799_1180# SG_DVDD SG_DVSS DOUT sky130_fd_pr__pfet_01v8_6QYSWZ
XXM8 SG_DVDD m1_3800_300# DOUT SG_DVSS sky130_fd_pr__nfet_01v8_723X3M
XXC4 SG_DVSS SG_DVDD sky130_fd_pr__cap_mim_m3_1_MPZGNS
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_JULQJE a_n287_n3288# a_n345_n3200# a_187_n3288#
+ a_n187_n3200# a_129_n3200# a_29_n3288# a_287_n3200# a_n129_n3288# a_n29_n3200# a_n479_n3422#
X0 a_287_n3200# a_187_n3288# a_129_n3200# a_n479_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=9.28 pd=64.58 as=4.64 ps=32.29 w=32 l=0.5
X1 a_n29_n3200# a_n129_n3288# a_n187_n3200# a_n479_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X2 a_n187_n3200# a_n287_n3288# a_n345_n3200# a_n479_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=9.28 ps=64.58 w=32 l=0.5
X3 a_129_n3200# a_29_n3288# a_n29_n3200# a_n479_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_844AHT a_n1135_n3200# a_1135_n3288# a_n445_n3288#
+ a_n919_n3288# a_n1551_n3288# a_n503_n3200# a_n1609_n3200# a_1609_n3288# a_819_n3288#
+ a_345_n3288# a_n287_n3288# a_n1393_n3288# a_n1867_n3288# a_2025_n3200# a_n345_n3200#
+ a_n819_n3200# a_n1451_n3200# a_1451_n3288# a_187_n3288# a_n761_n3288# a_n1925_n3200#
+ a_1925_n3288# a_n187_n3200# a_1293_n3288# a_661_n3288# a_n1293_n3200# a_n1767_n3200#
+ a_1767_n3288# a_2341_n3200# a_n661_n3200# a_977_n3288# a_n2025_n3288# a_2183_n3200#
+ a_n977_n3200# a_2499_n3200# a_n2341_n3288# a_n2183_n3288# a_n2691_n3422# a_n2241_n3200#
+ a_2241_n3288# a_n2499_n3288# a_n2083_n3200# a_2083_n3288# a_n2557_n3200# a_129_n3200#
+ a_29_n3288# a_n2399_n3200# a_2399_n3288# a_603_n3200# a_1709_n3200# a_1235_n3200#
+ a_919_n3200# a_445_n3200# a_1077_n3200# a_1551_n3200# a_287_n3200# a_n129_n3288#
+ a_n1235_n3288# a_761_n3200# a_n29_n3200# a_n603_n3288# a_n1709_n3288# a_1867_n3200#
+ a_1393_n3200# a_503_n3288# a_n1077_n3288#
X0 a_761_n3200# a_661_n3288# a_603_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X1 a_1867_n3200# a_1767_n3288# a_1709_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X2 a_2499_n3200# a_2399_n3288# a_2341_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=9.28 pd=64.58 as=4.64 ps=32.29 w=32 l=0.5
X3 a_n2241_n3200# a_n2341_n3288# a_n2399_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X4 a_n503_n3200# a_n603_n3288# a_n661_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X5 a_287_n3200# a_187_n3288# a_129_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X6 a_n661_n3200# a_n761_n3288# a_n819_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X7 a_n1135_n3200# a_n1235_n3288# a_n1293_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X8 a_n1293_n3200# a_n1393_n3288# a_n1451_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X9 a_n1609_n3200# a_n1709_n3288# a_n1767_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X10 a_n29_n3200# a_n129_n3288# a_n187_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X11 a_1551_n3200# a_1451_n3288# a_1393_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X12 a_2183_n3200# a_2083_n3288# a_2025_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X13 a_n2399_n3200# a_n2499_n3288# a_n2557_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=9.28 ps=64.58 w=32 l=0.5
X14 a_n1767_n3200# a_n1867_n3288# a_n1925_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X15 a_n187_n3200# a_n287_n3288# a_n345_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X16 a_2025_n3200# a_1925_n3288# a_1867_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X17 a_129_n3200# a_29_n3288# a_n29_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X18 a_445_n3200# a_345_n3288# a_287_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X19 a_919_n3200# a_819_n3288# a_761_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X20 a_n1925_n3200# a_n2025_n3288# a_n2083_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X21 a_n2083_n3200# a_n2183_n3288# a_n2241_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X22 a_n1451_n3200# a_n1551_n3288# a_n1609_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X23 a_1077_n3200# a_977_n3288# a_919_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X24 a_2341_n3200# a_2241_n3288# a_2183_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X25 a_n345_n3200# a_n445_n3288# a_n503_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X26 a_n819_n3200# a_n919_n3288# a_n977_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X27 a_n977_n3200# a_n1077_n3288# a_n1135_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X28 a_1235_n3200# a_1135_n3288# a_1077_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X29 a_603_n3200# a_503_n3288# a_445_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X30 a_1393_n3200# a_1293_n3288# a_1235_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X31 a_1709_n3200# a_1609_n3288# a_1551_n3200# a_n2691_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_KDBUUD a_50_n3200# a_n242_n3422# a_n50_n3288#
+ a_n108_n3200#
X0 a_50_n3200# a_n50_n3288# a_n108_n3200# a_n242_n3422# sky130_fd_pr__nfet_g5v0d10v5 ad=9.28 pd=64.58 as=9.28 ps=64.58 w=32 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YNEQJ5 a_50_n800# a_n108_n800# a_n50_n888# a_n242_n1022#
X0 a_50_n800# a_n50_n888# a_n108_n800# a_n242_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3 a_n242_n622# a_50_n400# a_n108_n400# a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n242_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH a_n345_n3200# a_29_n3297# a_n187_n3200#
+ a_n129_n3297# a_n287_n3297# a_187_n3297# w_n545_n3497# a_129_n3200# a_287_n3200#
+ a_n29_n3200#
X0 a_287_n3200# a_187_n3297# a_129_n3200# w_n545_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=9.28 pd=64.58 as=4.64 ps=32.29 w=32 l=0.5
X1 a_n29_n3200# a_n129_n3297# a_n187_n3200# w_n545_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X2 a_n187_n3200# a_n287_n3297# a_n345_n3200# w_n545_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=9.28 ps=64.58 w=32 l=0.5
X3 a_129_n3200# a_29_n3297# a_n29_n3200# w_n545_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_86VAEW a_n35_n1132# a_n189_n1286# a_n35_700#
X0 a_n35_700# a_n35_n1132# a_n189_n1286# sky130_fd_pr__res_xhigh_po_0p35 l=7.16
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_NH48NT a_n189_n866# a_n35_n712# a_n35_280#
X0 a_n35_280# a_n35_n712# a_n189_n866# sky130_fd_pr__res_xhigh_po_0p35 l=2.96
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQSVLT a_n1135_n3200# a_n2183_n3297# a_n503_n3200#
+ a_n1609_n3200# a_2241_n3297# a_n2499_n3297# a_2083_n3297# a_2025_n3200# a_n345_n3200#
+ a_n819_n3200# a_n1451_n3200# a_n1925_n3200# a_29_n3297# w_n2757_n3497# a_n187_n3200#
+ a_2399_n3297# a_n1293_n3200# a_n1767_n3200# a_2341_n3200# a_n661_n3200# a_2183_n3200#
+ a_n977_n3200# a_n129_n3297# a_2499_n3200# a_n1235_n3297# a_n1709_n3297# a_n603_n3297#
+ a_n1077_n3297# a_503_n3297# a_n445_n3297# a_n2241_n3200# a_1609_n3297# a_1135_n3297#
+ a_n919_n3297# a_n1551_n3297# a_345_n3297# a_n287_n3297# a_n2083_n3200# a_819_n3297#
+ a_n1393_n3297# a_n2557_n3200# a_187_n3297# a_n761_n3297# a_n1867_n3297# a_129_n3200#
+ a_1925_n3297# a_1451_n3297# a_n2399_n3200# a_661_n3297# a_603_n3200# a_1767_n3297#
+ a_1293_n3297# a_1709_n3200# a_1235_n3200# a_919_n3200# a_445_n3200# a_977_n3297#
+ a_n2025_n3297# a_1077_n3200# a_1551_n3200# a_287_n3200# a_761_n3200# a_n29_n3200#
+ a_n2341_n3297# a_1867_n3200# a_1393_n3200#
X0 a_761_n3200# a_661_n3297# a_603_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X1 a_1867_n3200# a_1767_n3297# a_1709_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X2 a_2499_n3200# a_2399_n3297# a_2341_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=9.28 pd=64.58 as=4.64 ps=32.29 w=32 l=0.5
X3 a_n2241_n3200# a_n2341_n3297# a_n2399_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X4 a_n503_n3200# a_n603_n3297# a_n661_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X5 a_287_n3200# a_187_n3297# a_129_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X6 a_n661_n3200# a_n761_n3297# a_n819_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X7 a_n1135_n3200# a_n1235_n3297# a_n1293_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X8 a_n1293_n3200# a_n1393_n3297# a_n1451_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X9 a_n1609_n3200# a_n1709_n3297# a_n1767_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X10 a_n29_n3200# a_n129_n3297# a_n187_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X11 a_1551_n3200# a_1451_n3297# a_1393_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X12 a_2183_n3200# a_2083_n3297# a_2025_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X13 a_n187_n3200# a_n287_n3297# a_n345_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X14 a_n2399_n3200# a_n2499_n3297# a_n2557_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=9.28 ps=64.58 w=32 l=0.5
X15 a_n1767_n3200# a_n1867_n3297# a_n1925_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X16 a_2025_n3200# a_1925_n3297# a_1867_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X17 a_129_n3200# a_29_n3297# a_n29_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X18 a_445_n3200# a_345_n3297# a_287_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X19 a_919_n3200# a_819_n3297# a_761_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X20 a_n1925_n3200# a_n2025_n3297# a_n2083_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X21 a_n2083_n3200# a_n2183_n3297# a_n2241_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X22 a_n1451_n3200# a_n1551_n3297# a_n1609_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X23 a_1077_n3200# a_977_n3297# a_919_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X24 a_2341_n3200# a_2241_n3297# a_2183_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X25 a_n345_n3200# a_n445_n3297# a_n503_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X26 a_n819_n3200# a_n919_n3297# a_n977_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X27 a_n977_n3200# a_n1077_n3297# a_n1135_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X28 a_1235_n3200# a_1135_n3297# a_1077_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X29 a_603_n3200# a_503_n3297# a_445_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X30 a_1393_n3200# a_1293_n3297# a_1235_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
X31 a_1709_n3200# a_1609_n3297# a_1551_n3200# w_n2757_n3497# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.29 as=4.64 ps=32.29 w=32 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCTT89 m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt vittoz_pierce_osc XOUT SG_AVDD EG_AVDD XIN EG_IBIAS AOUT SG_AVSS EG_AVSS
XXM12 m1_360_280# m1_n30_n90# m1_360_280# EG_AVSS EG_AVSS m1_360_280# m1_n30_n90#
+ m1_360_280# m1_n30_n90# EG_AVSS sky130_fd_pr__nfet_g5v0d10v5_JULQJE
XXM14 m1_2803_2950# m1_360_280# m1_360_280# m1_360_280# m1_360_280# m1_2803_2950#
+ m1_1740_7710# m1_360_280# m1_360_280# m1_360_280# m1_360_280# m1_360_280# m1_360_280#
+ m1_2803_2950# m1_1740_7710# m1_2803_2950# m1_2803_2950# m1_360_280# m1_360_280#
+ m1_360_280# m1_1740_7710# m1_360_280# m1_2803_2950# m1_360_280# m1_360_280# m1_1740_7710#
+ m1_2803_2950# m1_360_280# m1_2803_2950# m1_1740_7710# m1_360_280# m1_360_280# m1_1740_7710#
+ m1_1740_7710# m1_1740_7710# m1_360_280# m1_360_280# EG_AVSS m1_1740_7710# m1_360_280#
+ m1_360_280# m1_2803_2950# m1_360_280# m1_1740_7710# m1_2803_2950# m1_360_280# m1_2803_2950#
+ m1_360_280# m1_1740_7710# m1_2803_2950# m1_1740_7710# m1_1740_7710# m1_2803_2950#
+ m1_2803_2950# m1_1740_7710# m1_1740_7710# m1_360_280# m1_360_280# m1_2803_2950#
+ m1_1740_7710# m1_360_280# m1_360_280# m1_1740_7710# m1_2803_2950# m1_360_280# m1_360_280#
+ sky130_fd_pr__nfet_g5v0d10v5_844AHT
XXM13 EG_AVSS EG_AVSS XIN XOUT sky130_fd_pr__nfet_g5v0d10v5_KDBUUD
XXM15 EG_IBIAS m1_2803_2950# EG_IBIAS EG_AVSS EG_AVSS EG_IBIAS m1_2803_2950# EG_IBIAS
+ m1_2803_2950# EG_AVSS sky130_fd_pr__nfet_g5v0d10v5_JULQJE
XXM16 EG_AVSS EG_IBIAS EG_IBIAS EG_AVSS sky130_fd_pr__nfet_g5v0d10v5_YNEQJ5
XXM17 SG_AVSS SG_AVSS AOUT XIN sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3
XXM18 SG_AVDD m1_1740_7710# AOUT m1_1740_7710# m1_1740_7710# m1_1740_7710# SG_AVDD
+ AOUT SG_AVDD SG_AVDD sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH
XXR1 m1_360_280# EG_AVSS m1_n30_n90# sky130_fd_pr__res_xhigh_po_0p35_86VAEW
XXR3 EG_AVSS XIN XOUT sky130_fd_pr__res_xhigh_po_0p35_NH48NT
XXM9 XOUT m1_1740_7710# XOUT EG_AVDD m1_1740_7710# m1_1740_7710# m1_1740_7710# XOUT
+ EG_AVDD XOUT XOUT EG_AVDD m1_1740_7710# EG_AVDD XOUT m1_1740_7710# EG_AVDD XOUT
+ XOUT EG_AVDD EG_AVDD EG_AVDD m1_1740_7710# EG_AVDD m1_1740_7710# m1_1740_7710# m1_1740_7710#
+ m1_1740_7710# m1_1740_7710# m1_1740_7710# EG_AVDD m1_1740_7710# m1_1740_7710# m1_1740_7710#
+ m1_1740_7710# m1_1740_7710# m1_1740_7710# XOUT m1_1740_7710# m1_1740_7710# EG_AVDD
+ m1_1740_7710# m1_1740_7710# m1_1740_7710# XOUT m1_1740_7710# m1_1740_7710# XOUT
+ m1_1740_7710# EG_AVDD m1_1740_7710# m1_1740_7710# XOUT EG_AVDD EG_AVDD XOUT m1_1740_7710#
+ m1_1740_7710# XOUT EG_AVDD EG_AVDD XOUT EG_AVDD m1_1740_7710# EG_AVDD XOUT sky130_fd_pr__pfet_g5v0d10v5_AQSVLT
XXC1 EG_AVSS m1_n30_n90# sky130_fd_pr__cap_mim_m3_1_VCTT89
XXC2 m1_360_280# XIN sky130_fd_pr__cap_mim_m3_1_MPZGNS
XXC3 EG_AVSS EG_AVDD sky130_fd_pr__cap_mim_m3_1_MPZGNS
XXC4 SG_AVSS SG_AVDD sky130_fd_pr__cap_mim_m3_1_MPZGNS
XXC7 EG_AVSS m1_360_280# sky130_fd_pr__cap_mim_m3_1_MPZGNS
XXC8 SG_AVSS AOUT sky130_fd_pr__cap_mim_m3_1_VCTT89
XXM10 EG_AVDD m1_1740_7710# m1_n30_n90# m1_1740_7710# m1_1740_7710# m1_1740_7710#
+ EG_AVDD m1_n30_n90# EG_AVDD EG_AVDD sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH
XXM11 EG_AVDD m1_1740_7710# m1_1740_7710# m1_1740_7710# m1_1740_7710# m1_1740_7710#
+ EG_AVDD m1_1740_7710# EG_AVDD EG_AVDD sky130_fd_pr__pfet_g5v0d10v5_E4ZTVH
.ends

.subckt sky130_ht_ip__hsxo_cpz1 XOUT XIN ENA STDBY DOUT AVDD DVDD DVSS IBIAS power_gating_0/EG_AVSS
+ AVSS GUARD power_gating_0/SG_AVSS
Xpower_gating_0 DOUT power_gating_0/SG_AVDD power_gating_0/EG_IBIAS power_gating_0/SG_DVDD
+ AVDD power_gating_0/EG_AVDD ENA GUARD power_gating_0/SG_AVSS STDBY power_gating_0/EG_AVSS
+ XIN GUARD AVSS DVDD IBIAS DVSS power_gating
Xschmitt_trigger_pullmid_0 power_gating_0/SG_DVDD schmitt_trigger_pullmid_0/AIN DOUT
+ GUARD schmitt_trigger_pullmid
Xsky130_fd_pr__cap_mim_m3_1_MPZGNS_0 schmitt_trigger_pullmid_0/AIN vittoz_pierce_osc_0/AOUT
+ sky130_fd_pr__cap_mim_m3_1_MPZGNS
Xvittoz_pierce_osc_0 XOUT power_gating_0/SG_AVDD power_gating_0/EG_AVDD XIN power_gating_0/EG_IBIAS
+ vittoz_pierce_osc_0/AOUT power_gating_0/SG_AVSS power_gating_0/EG_AVSS vittoz_pierce_osc
.ends

.subckt isolated_switch_ena1v8 on dvdd in out avdd dvss avss
Xsky130_fd_pr__diode_pw2nd_05v5_HTFGEA_0 dvss on sky130_fd_pr__diode_pw2nd_05v5_HTFGEA
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 on dvdd dvss dvss avdd avdd isolated_switch_0/on
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xisolated_switch_0 isolated_switch_0/on avss out in avdd isolated_switch
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_LV9PDH a_8742_125# a_n3732_n557# a_1560_125#
+ a_3828_n557# a_n7512_n557# a_804_n557# a_7608_n557# a_n4110_n557# a_3072_125# a_4206_n557#
+ a_4584_125# a_n4110_125# a_6096_125# a_n5622_125# a_6852_n557# a_n4866_n557# a_n1464_n557#
+ a_3450_n557# a_48_125# a_n8646_n557# a_7230_n557# a_n5244_n557# a_n7134_125# a_n8646_125#
+ a_n1464_125# a_n9024_n557# a_n2976_125# a_804_125# a_2316_125# a_3828_125# a_n7890_n557#
+ a_5340_125# a_7986_n557# a_n4488_125# a_4584_n557# a_n2598_n557# a_1182_n557# a_6852_125#
+ a_8364_n557# a_n6378_n557# a_8364_125# a_1182_125# a_2694_125# a_n2220_125# a_n1842_n557#
+ a_48_n557# a_1938_n557# a_n3732_125# a_n708_125# a_n5622_n557# a_n2220_n557# a_5718_n557#
+ a_2316_n557# a_6096_n557# a_n5244_125# a_n6000_n557# a_n6756_125# a_7608_125# a_n8268_125#
+ a_n2976_n557# a_4962_n557# a_n1086_125# a_1560_n557# a_1938_125# a_n2598_125# a_3450_125#
+ a_4962_125# a_8742_n557# a_5340_n557# a_n6756_n557# a_426_125# a_n3354_n557# a_6474_125#
+ a_n7134_n557# a_426_n557# a_7986_125# a_n708_n557# a_n6000_125# a_n7512_125# a_2694_n557#
+ a_n1842_125# a_6474_n557# a_3072_n557# a_n4488_n557# a_n1086_n557# a_n330_125# a_n9024_125#
+ a_n3354_125# a_n8268_n557# a_n4866_125# a_n330_n557# a_n7890_125# a_4206_125# a_5718_125#
+ a_7230_125# VSUBS a_n6378_125#
X0 a_n8646_125# a_n8646_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X1 a_n6000_125# a_n6000_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X2 a_n1464_125# a_n1464_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X3 a_6474_125# a_6474_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X4 a_804_125# a_804_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X5 a_n7134_125# a_n7134_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X6 a_n4488_125# a_n4488_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X7 a_5718_125# a_5718_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X8 a_n1842_125# a_n1842_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X9 a_6852_125# a_6852_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X10 a_n7512_125# a_n7512_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X11 a_n4866_125# a_n4866_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X12 a_4206_125# a_4206_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X13 a_5340_125# a_5340_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X14 a_n330_125# a_n330_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X15 a_2694_125# a_2694_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X16 a_n7890_125# a_n7890_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X17 a_n3354_125# a_n3354_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X18 a_n2220_125# a_n2220_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X19 a_8364_125# a_8364_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X20 a_1182_125# a_1182_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X21 a_1938_125# a_1938_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X22 a_n9024_125# a_n9024_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X23 a_n708_125# a_n708_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X24 a_48_125# a_48_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X25 a_n6378_125# a_n6378_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X26 a_n3732_125# a_n3732_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X27 a_7608_125# a_7608_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X28 a_8742_125# a_8742_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X29 a_1560_125# a_1560_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X30 a_n6756_125# a_n6756_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X31 a_7230_125# a_7230_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X32 a_4584_125# a_4584_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X33 a_n5244_125# a_n5244_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X34 a_n4110_125# a_n4110_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X35 a_n2598_125# a_n2598_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X36 a_3072_125# a_3072_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X37 a_3828_125# a_3828_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X38 a_4962_125# a_4962_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X39 a_n8268_125# a_n8268_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X40 a_n5622_125# a_n5622_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X41 a_n2976_125# a_n2976_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X42 a_n1086_125# a_n1086_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X43 a_6096_125# a_6096_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X44 a_7986_125# a_7986_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X45 a_426_125# a_426_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X46 a_2316_125# a_2316_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X47 a_3450_125# a_3450_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_H3F4MM a_1182_1930# a_n4488_n1826# a_7986_n1826#
+ a_n6378_n2362# a_n7890_5150# a_n7890_n5582# a_7986_5150# a_4584_5150# a_n2598_5150#
+ a_1182_5150# a_8364_1930# a_n6378_1930# a_n4866_n1826# a_n6756_n2362# a_8364_5150#
+ a_n6378_5150# a_n2598_n1826# a_n6000_n5582# a_n4488_n2362# a_n3732_1394# a_7986_n2362#
+ a_3828_1394# a_426_n5582# a_7230_n5582# a_7608_n5582# a_n2976_n1826# a_n4866_n2362#
+ a_n7512_1394# a_n4110_1394# a_804_1394# a_7608_1394# a_4206_1394# a_4206_n1826#
+ a_n1842_1930# a_n4110_n5582# a_804_n5582# a_n2598_n2362# a_48_1930# a_1938_1930#
+ a_5340_n5582# a_n1842_5150# a_5718_n5582# a_48_5150# a_1938_5150# a_n5622_1930#
+ a_n2976_n2362# a_n2220_1930# a_5718_1930# a_3072_n5582# a_2316_1930# a_n9024_n1826#
+ a_6096_1930# a_2316_n1826# a_4206_n2362# a_n2220_n5582# a_n5622_5150# a_n2220_5150#
+ a_5718_5150# a_2316_5150# a_6852_1394# a_n6000_1930# a_6096_5150# a_n4866_1394#
+ a_3450_1394# a_3450_n5582# a_3828_n5582# a_n1464_1394# a_n8268_n5582# a_n6000_5150#
+ a_1182_n5582# a_n7134_n1826# a_n9024_n2362# a_2316_n2362# a_n8646_1394# a_7230_1394#
+ a_n5244_1394# a_8364_n1826# a_4962_1930# a_n2976_1930# a_1560_1930# a_n8646_n5582#
+ a_1560_n5582# a_n7512_n1826# a_1938_n5582# a_6096_n1826# a_n9024_1394# a_4962_5150#
+ a_n2976_5150# a_n6378_n5582# a_n5244_n1826# a_n7134_n2362# a_1560_5150# a_8742_n1826#
+ a_8742_1930# a_n6756_1930# a_5340_1930# a_n3354_1930# a_n330_n1826# a_6474_n1826#
+ a_n708_n1826# a_8364_n2362# a_8742_5150# a_n6756_n5582# a_n6756_5150# a_n5622_n1826#
+ a_5340_5150# a_n7512_n2362# a_48_n1826# a_n7890_1394# a_n3354_5150# a_6096_n2362#
+ a_n7134_1930# a_7986_1394# a_n4488_n5582# a_426_1930# a_4584_1394# a_7986_n5582#
+ a_n3354_n1826# a_n2598_1394# a_6852_n1826# a_n5244_n2362# a_8742_n2362# a_1182_1394#
+ a_n708_1930# a_n7134_5150# a_n1086_n1826# a_426_5150# a_4584_n1826# a_n330_n2362#
+ a_6474_n2362# a_n708_n2362# a_8364_1394# a_n4866_n5582# a_n3732_n1826# a_n6378_1394#
+ a_n5622_n2362# a_48_n2362# a_n708_5150# a_2694_1930# a_n2598_n5582# a_n1464_n1826#
+ a_4962_n1826# a_n3354_n2362# a_6852_n2362# a_2694_5150# a_2694_n1826# a_n1086_n2362#
+ a_4584_n2362# a_6474_1930# a_n2976_n5582# a_n4488_1930# a_n1842_n1826# a_n3732_n2362#
+ a_3072_1930# a_n1086_1930# a_4206_n5582# a_6474_5150# a_n1464_n2362# a_4962_n2362#
+ a_n4488_5150# a_3072_5150# a_n1842_1394# a_n1086_5150# a_n8268_1930# a_48_1394#
+ a_1938_1394# a_2694_n2362# a_n330_1930# a_n1842_n2362# a_n8268_5150# a_n5622_1394#
+ a_n9024_n5582# a_n2220_1394# a_2316_n5582# a_5718_1394# a_n7890_n1826# a_n330_5150#
+ a_2316_1394# a_6096_1394# a_n6000_1394# a_n3732_1930# a_n7134_n5582# a_3828_1930#
+ a_n6000_n1826# a_n7890_n2362# a_n3732_5150# a_8364_n5582# a_426_n1826# a_7230_n1826#
+ a_3828_5150# a_7608_n1826# a_n7512_1930# a_n7512_n5582# a_n4110_1930# a_804_1930#
+ a_7608_1930# a_4962_1394# a_n2976_1394# a_4206_1930# a_1560_1394# a_6096_n5582#
+ a_n7512_5150# a_n5244_n5582# a_n4110_n1826# a_8742_n5582# a_804_n1826# a_n6000_n2362#
+ a_n4110_5150# a_804_5150# a_7608_5150# a_4206_5150# a_8742_1394# a_n6756_1394# a_5340_1394#
+ a_n3354_1394# a_6474_n5582# a_n330_n5582# a_n708_n5582# a_5340_n1826# a_426_n2362#
+ a_5718_n1826# a_7230_n2362# a_7608_n2362# a_n5622_n5582# a_48_n5582# a_3072_n1826#
+ a_n7134_1394# a_n3354_n5582# a_6852_n5582# a_n2220_n1826# a_n4110_n2362# a_804_n2362#
+ a_426_1394# a_6852_1930# a_n4866_1930# a_3450_1930# a_n1464_1930# a_n1086_n5582#
+ a_4584_n5582# a_n708_1394# a_3450_n1826# a_5340_n2362# a_3828_n1826# a_5718_n2362#
+ a_n3732_n5582# a_6852_5150# a_n4866_5150# a_3450_5150# a_n1464_5150# a_n8268_n1826#
+ a_1182_n1826# a_n8646_1930# a_3072_n2362# a_7230_1930# a_n5244_1930# a_n1464_n5582#
+ a_4962_n5582# a_n2220_n2362# a_2694_1394# a_n8646_5150# a_7230_5150# a_2694_n5582#
+ a_n8646_n1826# a_n5244_5150# a_1560_n1826# a_1938_n1826# a_3450_n2362# a_3828_n2362#
+ a_n9024_1930# a_n1842_n5582# a_6474_1394# a_n4488_1394# a_3072_1394# a_n6378_n1826#
+ a_n8268_n2362# a_n1086_1394# a_1182_n2362# a_n9024_5150# a_n8268_1394# a_n7890_1930#
+ a_n6756_n1826# a_n8646_n2362# a_1560_n2362# a_1938_n2362# a_7986_1930# VSUBS a_4584_1930#
+ a_n2598_1930# a_n330_1394#
X0 a_n1464_n2362# a_n1464_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X1 a_n3732_n2362# a_n3732_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X2 a_426_n2362# a_426_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X3 a_n4110_5150# a_n4110_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X4 a_n5244_5150# a_n5244_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X5 a_n2598_5150# a_n2598_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X6 a_3072_5150# a_3072_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X7 a_3828_5150# a_3828_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X8 a_4962_5150# a_4962_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X9 a_n9024_1394# a_n9024_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X10 a_6474_1394# a_6474_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X11 a_n8268_5150# a_n8268_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X12 a_8742_1394# a_8742_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X13 a_5718_1394# a_5718_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X14 a_n330_1394# a_n330_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X15 a_n9024_n2362# a_n9024_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X16 a_3072_1394# a_3072_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X17 a_n7890_1394# a_n7890_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X18 a_n5622_5150# a_n5622_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X19 a_5340_1394# a_5340_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X20 a_2316_1394# a_2316_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X21 a_n1086_5150# a_n1086_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X22 a_6096_5150# a_6096_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X23 a_6474_n2362# a_6474_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X24 a_8742_n2362# a_8742_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X25 a_5718_n2362# a_5718_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X26 a_n330_n2362# a_n330_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X27 a_7986_5150# a_7986_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X28 a_n4488_1394# a_n4488_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X29 a_n2976_5150# a_n2976_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X30 a_2316_5150# a_2316_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X31 a_n6756_1394# a_n6756_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X32 a_426_5150# a_426_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X33 a_3450_5150# a_3450_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X34 a_3072_n2362# a_3072_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X35 a_n7890_n2362# a_n7890_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X36 a_5340_n2362# a_5340_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X37 a_2316_n2362# a_2316_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X38 a_n1086_1394# a_n1086_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X39 a_n3354_1394# a_n3354_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X40 a_n4488_n2362# a_n4488_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X41 a_n5622_1394# a_n5622_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X42 a_n6756_n2362# a_n6756_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X43 a_n1086_n2362# a_n1086_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X44 a_n8646_5150# a_n8646_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X45 a_n3354_n2362# a_n3354_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X46 a_n5622_n2362# a_n5622_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X47 a_n6000_5150# a_n6000_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X48 a_6474_5150# a_6474_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X49 a_n1464_5150# a_n1464_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X50 a_804_5150# a_804_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X51 a_n7134_5150# a_n7134_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X52 a_6096_1394# a_6096_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X53 a_n4488_5150# a_n4488_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X54 a_8364_1394# a_8364_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X55 a_7608_1394# a_7608_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X56 a_n1842_5150# a_n1842_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X57 a_5718_5150# a_5718_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X58 a_6852_5150# a_6852_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X59 a_6096_n2362# a_6096_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X60 a_7230_1394# a_7230_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X61 a_4206_1394# a_4206_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X62 a_8364_n2362# a_8364_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X63 a_7608_n2362# a_7608_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X64 a_n6378_1394# a_n6378_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X65 a_n8646_1394# a_n8646_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X66 a_7230_n2362# a_7230_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X67 a_4206_n2362# a_4206_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X68 a_n2220_1394# a_n2220_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X69 a_n5244_1394# a_n5244_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X70 a_n6378_n2362# a_n6378_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X71 a_n7512_1394# a_n7512_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X72 a_n7512_5150# a_n7512_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X73 a_n8646_n2362# a_n8646_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X74 a_2694_1394# a_2694_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X75 a_n4866_5150# a_n4866_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X76 a_4206_5150# a_4206_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X77 a_4962_1394# a_4962_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X78 a_1938_1394# a_1938_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X79 a_5340_5150# a_5340_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X80 a_n2220_n2362# a_n2220_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X81 a_n5244_n2362# a_n5244_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X82 a_n7512_n2362# a_n7512_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X83 a_n330_5150# a_n330_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X84 a_2694_5150# a_2694_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X85 a_1560_1394# a_1560_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X86 a_2694_n2362# a_2694_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X87 a_4962_n2362# a_4962_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X88 a_1938_n2362# a_1938_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X89 a_48_1394# a_48_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X90 a_n2976_1394# a_n2976_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X91 a_1560_n2362# a_1560_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X92 a_48_n2362# a_48_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X93 a_n7890_5150# a_n7890_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X94 a_n1842_1394# a_n1842_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X95 a_n2220_5150# a_n2220_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X96 a_n2976_n2362# a_n2976_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X97 a_n3354_5150# a_n3354_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X98 a_8364_5150# a_8364_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X99 a_804_1394# a_804_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X100 a_1182_5150# a_1182_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X101 a_n1842_n2362# a_n1842_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X102 a_1938_5150# a_1938_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X103 a_804_n2362# a_804_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X104 a_n708_5150# a_n708_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X105 a_48_5150# a_48_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X106 a_n9024_5150# a_n9024_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X107 a_n8268_1394# a_n8268_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X108 a_n6378_5150# a_n6378_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X109 a_n3732_5150# a_n3732_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X110 a_7608_5150# a_7608_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X111 a_8742_5150# a_8742_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X112 a_7986_1394# a_7986_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X113 a_n4110_1394# a_n4110_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X114 a_n7134_1394# a_n7134_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X115 a_n8268_n2362# a_n8268_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X116 a_4584_1394# a_4584_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X117 a_1560_5150# a_1560_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X118 a_6852_1394# a_6852_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X119 a_3828_1394# a_3828_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X120 a_7986_n2362# a_7986_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X121 a_n4110_n2362# a_n4110_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X122 a_n7134_n2362# a_n7134_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X123 a_n708_1394# a_n708_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X124 a_1182_1394# a_1182_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X125 a_n6000_1394# a_n6000_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X126 a_3450_1394# a_3450_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X127 a_4584_n2362# a_4584_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X128 a_6852_n2362# a_6852_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X129 a_3828_n2362# a_3828_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X130 a_n2598_1394# a_n2598_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X131 a_n708_n2362# a_n708_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X132 a_n4866_1394# a_n4866_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X133 a_n6756_5150# a_n6756_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X134 a_1182_n2362# a_1182_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X135 a_n6000_n2362# a_n6000_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X136 a_7230_5150# a_7230_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X137 a_3450_n2362# a_3450_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X138 a_n1464_1394# a_n1464_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X139 a_4584_5150# a_4584_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X140 a_n2598_n2362# a_n2598_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X141 a_n3732_1394# a_n3732_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X142 a_n4866_n2362# a_n4866_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X143 a_426_1394# a_426_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8 a_300_n300# a_n492_n522# a_n358_n300#
+ a_n300_n388#
X0 a_300_n300# a_n300_n388# a_n358_n300# a_n492_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=3
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_F6RBXN a_n147_n172# a_n45_n70#
X0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
.ends

.subckt voltage_divider out_0000 out_0001 out_0010 out_0011 out_0100 out_0101 out_0110
+ out_0111 out_1000 out_1001 out_1010 out_1011 out_1100 out_1101 out_1110 out_1111
+ ena avdd avss
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_0 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_2 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_H3F4MM_0 m1_3399_9649# m1_7155_3979# m1_7155_16831#
+ m1_7155_2467# m1_179_955# m1_10911_577# m1_179_16831# m1_179_13051# m1_179_6247#
+ m1_179_10027# m1_3399_17209# m1_3399_2467# m1_7155_3979# m1_7155_2089# m1_179_16831#
+ m1_179_2467# m1_7155_6247# m1_10911_2845# out_1110 m1_3935_5113# m1_7155_16831#
+ m1_3935_12673# out_0011 m1_10911_15697# m1_10911_16453# m1_7155_5491# out_1110 m1_3399_1333#
+ m1_3935_4357# m1_3935_9649# m1_3935_16453# m1_3935_12673# m1_7155_13051# m1_3399_6625#
+ out_1101 out_0010 out_1000 m1_3399_8893# m1_3399_10405# m1_10911_14185# m1_179_7003#
+ m1_10911_14185# m1_179_8515# m1_179_10783# m1_3399_3223# out_1010 m1_3399_6625#
+ m1_3399_14185# m1_10911_11917# m1_3399_11161# avss m1_3399_14941# m1_7155_10783#
+ m1_7691_13051# out_0111 m1_179_3223# m1_179_6247# m1_179_14563# m1_179_10783# m1_3935_15697#
+ m1_3399_2845# m1_179_14563# m1_3399_3979# m1_3935_11917# m1_10911_11917# m1_10911_12673#
+ m1_3935_7381# m1_10911_577# m1_179_2467# out_0010 m1_7155_1711# avss m1_7691_10783#
+ m1_3399_199# m1_3935_15697# m1_3399_3601# m1_7155_17209# m1_3399_13429# m1_3399_5869#
+ m1_3399_10405# m1_10901_199# out_0001 m1_7155_1333# out_0001 m1_7155_14563# avss
+ m1_179_13807# m1_179_5491# m1_10911_2089# m1_7155_3601# m1_7155_1711# m1_179_10027#
+ avss avss m1_3399_2089# m1_3399_14185# m1_3399_5113# m1_7155_8515# m1_7155_15319#
+ m1_7155_7759# m1_7155_17209# avss m1_10911_2089# m1_179_1711# m1_7155_3223# m1_179_13807#
+ m1_7155_1333# m1_7155_8515# m1_3399_955# m1_179_5491# m1_7691_14563# m1_3399_1711#
+ m1_3935_16453# out_1101 m1_3399_8893# m1_3935_13429# m1_10911_16453# m1_7155_5491#
+ m1_3935_5869# m1_7155_15319# m1_7155_3601# avss m1_3935_9649# m1_3399_8137# m1_179_1711#
+ m1_7155_7759# m1_179_9271# m1_7155_13051# out_0100 m1_7691_15319# out_0101 m1_3399_17209#
+ out_1111 m1_7155_4735# m1_3399_2467# m1_7155_3223# out_0100 m1_179_7759# m1_3399_11161#
+ out_1001 m1_7155_7003# m1_7155_13807# out_1010 m1_7691_15319# m1_179_11539# m1_7155_11539#
+ out_0101 m1_7691_13051# m1_3399_14941# out_1001 m1_3399_4357# m1_7155_7003# out_1100
+ m1_3399_11917# m1_3399_7381# m1_10911_12673# m1_179_15319# m1_7691_7003# m1_7691_13807#
+ m1_179_3979# m1_179_11539# m1_3935_6625# m1_179_7759# m1_3399_577# m1_3935_8893#
+ m1_3935_10405# 51 m1_3399_8137# m1_7691_7003# m1_179_199# m1_3399_3223# avss m1_3935_6625#
+ out_0000 m1_3935_14185# m1_7155_955# m1_179_8515# m1_3935_11161# m1_3935_14941#
+ m1_3399_2845# m1_3399_5113# m1_10911_1333# m1_3399_12673# m1_7155_2845# m1_7155_955#
+ m1_179_4735# avdd m1_7155_9271# m1_7155_16075# m1_179_12295# m1_7155_16075# m1_3399_1333#
+ m1_10911_1333# m1_3399_4357# m1_3399_9649# m1_3399_16453# m1_3935_13429# m1_3935_5869#
+ m1_3399_12673# m1_3935_10405# m1_10911_14941# m1_179_955# out_1111 m1_7155_4735#
+ avss m1_7155_9271# m1_7155_2845# m1_179_4735# m1_179_9271# m1_179_16075# m1_179_13051#
+ avss m1_3399_2089# m1_3935_14185# m1_3935_5113# m1_10911_14941# m1_10901_8137# m1_10901_8137#
+ m1_7155_13807# m1_7691_9271# m1_7155_14563# m1_7691_16075# m1_7691_16075# m1_10911_2845#
+ out_0011 m1_7155_11539# m1_3399_1711# out_1011 m1_10911_15697# m1_7155_6247# out_1100
+ m1_7691_9271# m1_3935_8893# m1_3399_15697# m1_3399_3979# m1_3399_11917# m1_3399_7381#
+ out_0110 m1_10911_13429# m1_3935_8137# m1_7155_12295# m1_7691_13807# m1_7155_12295#
+ m1_7691_14563# out_1011 m1_179_15319# m1_179_3979# m1_179_12295# m1_179_7003# m1_7155_577#
+ m1_7155_10027# m1_3399_199# 51 m1_3399_15697# m1_3399_3601# out_0110 m1_10911_13429#
+ out_1000 m1_3935_11161# m1_179_199# m1_179_16075# out_0000 m1_7155_199# m1_179_3223#
+ m1_7155_10027# m1_7155_10783# m1_7691_12295# m1_7691_12295# avss out_0111 m1_3935_14941#
+ m1_3935_4357# m1_3935_11917# m1_7155_2467# m1_7155_577# m1_3935_7381# m1_7691_10027#
+ avss m1_3399_577# m1_3399_955# m1_7155_2089# m1_7155_199# m1_7691_10027# m1_7691_10783#
+ m1_3399_16453# avss m1_3399_13429# m1_3399_5869# m1_3935_8137# sky130_fd_pr__res_xhigh_po_1p41_H3F4MM
Xsky130_fd_pr__nfet_g5v0d10v5_SB5CJ8_0 avss avss m1_10901_199# ena sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CY564Z a_300_n100# a_n492_n322# a_n358_n100#
+ a_n300_n188#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n492_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt trans_gate_m in ena_b ena out avdd vss
Xsky130_fd_pr__pfet_g5v0d10v5_6H9SQ3_1 ena_b out avdd in sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3
Xsky130_fd_pr__nfet_g5v0d10v5_CY564Z_0 out vss in ena sky130_fd_pr__nfet_g5v0d10v5_CY564Z
.ends

.subckt multiplexer in_0000 in_0001 in_0010 in_0011 in_0100 in_0101 in_0110 in_0111
+ vtrip_3 vtrip_3_b vtrip_2 vtrip_1 out vtrip_1_b vtrip_0 vtrip_0_b in_1000 in_1001
+ in_1010 in_1011 in_1100 in_1101 in_1110 in_1111 vtrip_2_b vss avdd
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_3 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_2 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_4 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_5 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_6 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_7 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_8 vss vtrip_2_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_9 vss vtrip_2 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_31 trans_gate_m_31/in vtrip_1 vtrip_1_b trans_gate_m_20/in avdd vss
+ trans_gate_m
Xtrans_gate_m_20 trans_gate_m_20/in vtrip_2 vtrip_2_b trans_gate_m_33/in avdd vss
+ trans_gate_m
Xtrans_gate_m_0 in_0010 vtrip_0 vtrip_0_b trans_gate_m_29/in avdd vss trans_gate_m
Xtrans_gate_m_1 in_0011 vtrip_0_b vtrip_0 trans_gate_m_29/in avdd vss trans_gate_m
Xtrans_gate_m_32 trans_gate_m_32/in vtrip_2 vtrip_2_b trans_gate_m_34/in avdd vss
+ trans_gate_m
Xtrans_gate_m_10 in_1000 vtrip_0 vtrip_0_b trans_gate_m_23/in avdd vss trans_gate_m
Xtrans_gate_m_21 trans_gate_m_5/out vtrip_1_b vtrip_1 trans_gate_m_32/in avdd vss
+ trans_gate_m
Xtrans_gate_m_2 in_0110 vtrip_0 vtrip_0_b trans_gate_m_3/out avdd vss trans_gate_m
Xtrans_gate_m_33 trans_gate_m_33/in vtrip_3 vtrip_3_b out avdd vss trans_gate_m
Xtrans_gate_m_11 in_1001 vtrip_0_b vtrip_0 trans_gate_m_23/in avdd vss trans_gate_m
Xtrans_gate_m_3 in_0111 vtrip_0_b vtrip_0 trans_gate_m_3/out avdd vss trans_gate_m
Xtrans_gate_m_12 in_0101 vtrip_0_b vtrip_0 trans_gate_m_27/in avdd vss trans_gate_m
Xtrans_gate_m_34 trans_gate_m_34/in vtrip_3_b vtrip_3 out avdd vss trans_gate_m
Xtrans_gate_m_23 trans_gate_m_23/in vtrip_1 vtrip_1_b trans_gate_m_32/in avdd vss
+ trans_gate_m
Xtrans_gate_m_13 in_0100 vtrip_0 vtrip_0_b trans_gate_m_27/in avdd vss trans_gate_m
Xtrans_gate_m_4 in_1011 vtrip_0_b vtrip_0 trans_gate_m_5/out avdd vss trans_gate_m
Xtrans_gate_m_14 in_0001 vtrip_0_b vtrip_0 trans_gate_m_31/in avdd vss trans_gate_m
Xtrans_gate_m_25 trans_gate_m_3/out vtrip_1_b vtrip_1 trans_gate_m_28/in avdd vss
+ trans_gate_m
Xtrans_gate_m_5 in_1010 vtrip_0 vtrip_0_b trans_gate_m_5/out avdd vss trans_gate_m
Xtrans_gate_m_15 in_0000 vtrip_0 vtrip_0_b trans_gate_m_31/in avdd vss trans_gate_m
Xtrans_gate_m_27 trans_gate_m_27/in vtrip_1 vtrip_1_b trans_gate_m_28/in avdd vss
+ trans_gate_m
Xtrans_gate_m_37 trans_gate_m_37/in vtrip_2_b vtrip_2 trans_gate_m_34/in avdd vss
+ trans_gate_m
Xtrans_gate_m_6 in_1110 vtrip_0 vtrip_0_b trans_gate_m_7/out avdd vss trans_gate_m
Xtrans_gate_m_28 trans_gate_m_28/in vtrip_2_b vtrip_2 trans_gate_m_33/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_10 vss vtrip_3_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_7 in_1111 vtrip_0_b vtrip_0 trans_gate_m_7/out avdd vss trans_gate_m
Xtrans_gate_m_29 trans_gate_m_29/in vtrip_1_b vtrip_1 trans_gate_m_20/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_11 vss vtrip_3 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_18 trans_gate_m_9/out vtrip_1 vtrip_1_b trans_gate_m_37/in avdd vss
+ trans_gate_m
Xtrans_gate_m_8 in_1101 vtrip_0_b vtrip_0 trans_gate_m_9/out avdd vss trans_gate_m
Xtrans_gate_m_19 trans_gate_m_7/out vtrip_1_b vtrip_1 trans_gate_m_37/in avdd vss
+ trans_gate_m
Xtrans_gate_m_9 in_1100 vtrip_0 vtrip_0_b trans_gate_m_9/out avdd vss trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_1 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YHAZV5 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_37RBXE a_n147_n172# a_n45_n70#
X0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EEVBR7 a_n300_n288# a_300_n200# a_n492_n422#
+ a_n358_n200#
X0 a_300_n200# a_n300_n288# a_n358_n200# a_n492_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_MG6U6H a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9Q3 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt level_shifter in out out_b dvss avss M2 avdd
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0 out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1 out out_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__diode_pw2nd_05v5_37RBXE_0 dvss in sky130_fd_pr__diode_pw2nd_05v5_37RBXE
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0 in_b out avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1 in out_b avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_01v8_MG6U6H_0 dvss in_b in dvss sky130_fd_pr__nfet_01v8_MG6U6H
Xsky130_fd_pr__pfet_01v8_J2L9Q3_0 in in_b M2 M2 sky130_fd_pr__pfet_01v8_J2L9Q3
.ends

.subckt sky130_fd_pr__pfet_01v8_XTWSDC a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
.ends

.subckt sky130_fd_pr__nfet_01v8_7ZF23Z a_2000_n100# a_n2058_n100# a_n2000_n188# a_n2160_n274#
X0 a_2000_n100# a_n2000_n188# a_n2058_n100# a_n2160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_V433WY a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69BJMM a_n500_n188# a_500_n100# a_n692_n322#
+ a_n558_n100#
X0 a_500_n100# a_n500_n188# a_n558_n100# a_n692_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E7V9VM w_n758_n897# a_n558_n600# a_n500_n697#
+ a_500_n600#
X0 a_500_n600# a_n500_n697# a_n558_n600# w_n758_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=5
.ends

.subckt trans_gate in ena_b ena out vss avdd
XXM1 ena out vss in sky130_fd_pr__nfet_g5v0d10v5_69BJMM
XXM2 avdd out ena_b in sky130_fd_pr__pfet_g5v0d10v5_E7V9VM
.ends

.subckt sky130_fd_pr__pfet_01v8_C2YSV5 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9E5 w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_GGMWVD w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_CDT3CS a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
.ends

.subckt sky130_fd_pr__pfet_01v8_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397# a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_697RXD a_800_n100# a_n858_n100# a_n800_n188# a_n960_n274#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n960_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_4T6WVE a_100_n130# a_n292_n352# a_n158_n130#
+ a_n100_n218#
X0 a_100_n130# a_n100_n218# a_n158_n130# a_n292_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_6975WM a_800_n130# a_n992_n352# a_n858_n130#
+ a_n800_n218#
X0 a_800_n130# a_n800_n218# a_n858_n130# a_n992_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DEN7YK a_800_n100# a_n992_n322# a_n858_n100#
+ a_n800_n188#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n992_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_G3L97A w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_C8TQ3N a_n158_n300# a_n100_n388# a_n260_n474# a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n260_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt comp_hyst out vref vin ena ibias dvss dvdd
XXMD16[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM12 dvss net1 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
XXM14 dvss net2 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXM13 dvss net5 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
Xx1 ibias ena_b ena net5 dvss dvdd trans_gate
XXM15 ena net4 dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXM16 ena net3 dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXM17 dvss out ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXMD1[19] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM18 ena ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXMD1[18] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM19 dvss ena_b ena dvss sky130_fd_pr__nfet_01v8_V433WY
XXM6[3] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM3[1] dvdd net4 net4 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[17] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[2] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXM3[0] dvdd net4 net4 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[16] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[1] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM6[0] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXMD1[15] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[13] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[14] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[9] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[12] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[8] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[11] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[7] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[10] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[6] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XD1 dvss vref sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM7 dvdd net4 net2 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM9 dvdd dvdd net3 out sky130_fd_pr__pfet_01v8_3HBZVM
XXM8 dvss net2 net2 dvss sky130_fd_pr__nfet_01v8_697RXD
XXMDN13[7] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXM1[1] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXMD1[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM1[0] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM4[1] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMDN13[6] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMD1[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM4[0] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXMDN13[5] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[4] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN8[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMDN8[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMD16[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMD16[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[1] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[1] dvdd net4 net3 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[0] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[0] dvdd net4 net3 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMD8[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_G3L97A
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 dvss vin sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXM10 out net2 dvss dvss sky130_fd_pr__nfet_01v8_C8TQ3N
XXMD8[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_G3L97A
XXMD16[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM11 dvss net5 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
.ends

.subckt sky130_vbl_ip__overvoltage avdd dvdd ena vtrip[3] ibias vtrip[2] ovout vbg
+ vtrip[1] vtrip[0] dvss avss
Xvoltage_divider_0 multiplexer_0/in_0000 multiplexer_0/in_0001 multiplexer_0/in_0010
+ multiplexer_0/in_0011 multiplexer_0/in_0100 multiplexer_0/in_0101 multiplexer_0/in_0110
+ multiplexer_0/in_0111 multiplexer_0/in_1000 multiplexer_0/in_1001 multiplexer_0/in_1010
+ multiplexer_0/in_1011 multiplexer_0/in_1100 multiplexer_0/in_1101 multiplexer_0/in_1110
+ multiplexer_0/in_1111 ena avdd avss voltage_divider
Xmultiplexer_0 multiplexer_0/in_0000 multiplexer_0/in_0001 multiplexer_0/in_0010 multiplexer_0/in_0011
+ multiplexer_0/in_0100 multiplexer_0/in_0101 multiplexer_0/in_0110 multiplexer_0/in_0111
+ level_shifter_3/out level_shifter_3/out_b level_shifter_2/out level_shifter_1/out
+ vin level_shifter_1/out_b level_shifter_0/out level_shifter_0/out_b multiplexer_0/in_1000
+ multiplexer_0/in_1001 multiplexer_0/in_1010 multiplexer_0/in_1011 multiplexer_0/in_1100
+ multiplexer_0/in_1101 multiplexer_0/in_1110 multiplexer_0/in_1111 level_shifter_2/out_b
+ avss avdd multiplexer
Xlevel_shifter_0 vtrip[0] level_shifter_0/out level_shifter_0/out_b dvss avss dvdd
+ avdd level_shifter
Xlevel_shifter_1 vtrip[1] level_shifter_1/out level_shifter_1/out_b dvss avss dvdd
+ avdd level_shifter
Xlevel_shifter_2 vtrip[2] level_shifter_2/out level_shifter_2/out_b dvss avss dvdd
+ avdd level_shifter
Xlevel_shifter_3 vtrip[3] level_shifter_3/out level_shifter_3/out_b dvss avss dvdd
+ avdd level_shifter
Xcomp_hyst_0 ovout vbg vin ena ibias dvss dvdd comp_hyst
.ends

.subckt lvl_shift_invert in1v8 dvdd avdd outb3v3 out3v3 dvss
Xsky130_fd_sc_hvl__inv_2_0 out3v3 dvss dvss avdd avdd outb3v3 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 in1v8 dvdd dvss dvss avdd avdd out3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
.ends

.subckt sky130_fd_pr__nfet_01v8_QXBCRM a_n1000_n188# a_n1160_n274# a_1000_n100# a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B5H3CA w_n1196_n319# a_n1000_n197# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1196_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt buffer vdd input output vbias vss
XXM1 input vss m1_2942_n986# m1_772_n974# sky130_fd_pr__nfet_01v8_QXBCRM
XXM2 output vss output m1_2942_n986# sky130_fd_pr__nfet_01v8_QXBCRM
XXM3 vdd m1_772_n974# vdd m1_772_n974# sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM4 vdd m1_772_n974# output vdd sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM5 vbias vss m1_2942_n986# vss sky130_fd_pr__nfet_01v8_QXBCRM
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6VRZAW a_100_n536# w_n296_n1191# a_n100_675# a_100_336#
+ a_n158_n536# a_n158_772# a_n100_n633# a_n100_239# a_n100_n197# a_100_n100# a_n158_336#
+ a_100_n972# a_n158_n100# a_100_772# a_n158_n972# a_n100_n1069#
X0 a_100_336# a_n100_239# a_n158_336# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_772# a_n100_675# a_n158_772# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n536# a_n100_n633# a_n158_n536# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n972# a_n100_n1069# a_n158_n972# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_3VR9VM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_od_ip__tempsensor_ext_vp vbe2_out vbe1_out ena vbg vdd vss
Xx1 vdd x1/input vbe2_out ena vss buffer
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 vss vbg sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_1 vss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_2 vss vbe1_out sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xx2 vdd x2/input vbe1_out ena vss buffer
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_3 vss vbe2_out sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXQ_BR1 x1/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXQ_BL1 x2/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM22 vdd vdd m1_1668_n386# vdd x1/input x1/input m1_1668_n386# m1_1668_n386# m1_1668_n386#
+ vdd x1/input vdd x1/input vdd x1/input m1_1668_n386# sky130_fd_pr__pfet_01v8_lvt_6VRZAW
XXM11 vdd m1_1668_n386# vdd x2/input sky130_fd_pr__pfet_01v8_lvt_3VR9VM
XXM66 ena vss m1_772_n1144# vss sky130_fd_pr__nfet_01v8_QXBCRM
XXM88 vdd m1_420_n380# vdd m1_420_n380# sky130_fd_pr__pfet_01v8_3HMWVM
XXM77 vdd m1_420_n380# m1_1668_n386# vdd sky130_fd_pr__pfet_01v8_3HMWVM
XXM33 vdd ena m1_1668_n386# vdd sky130_fd_pr__pfet_01v8_3HMWVM
XXM55 vss m1_1668_n386# m1_772_n1144# m1_1668_n386# sky130_fd_pr__nfet_01v8_69TQ3K
XXM44 vss m1_772_n1144# m1_420_n380# vbg sky130_fd_pr__nfet_01v8_69TQ3K
.ends

.subckt bbp__M5 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bbp__M6 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bbp__M4 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bbp__M4_nc w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bb__pmirr vbn vbp ibp vdd
Xbbp__M5_2 vdd vbp vdd vbp bbp__M5
Xbbp__M5_3 vdd vdd vbp vbp bbp__M5
Xbbp__M5_4 vdd vbp vdd vbp bbp__M5
Xbbp__M5_5 vdd vdd vbp vbp bbp__M5
Xbbp__M5_6 vdd vbp vdd vbp bbp__M5
Xbbp__M5_7 vdd vdd vbp vbp bbp__M5
Xbbp__M6_0 vdd ibp vdd vbp bbp__M6
Xbbp__M6_1 vdd vdd ibp vbp bbp__M6
Xbbp__M4_0 vdd vbn vdd vbp bbp__M4
Xbbp__M4_1 vdd vdd vbn vbp bbp__M4
Xbbp__M4_3 vdd vbn vdd vbp bbp__M4
Xbbp__M4_2 vdd vdd vbn vbp bbp__M4
Xbbp__M4_nc_0 vdd vbn vdd vbp bbp__M4_nc
Xbbp__M4_nc_1 vdd vbn vdd vbp bbp__M4_nc
Xbbp__M4_nc_2 vdd vdd vbn vbp bbp__M4_nc
Xbbp__M4_nc_3 vdd vdd vbn vbp bbp__M4_nc
Xbbp__M5_0 vdd vbp vdd vbp bbp__M5
Xbbp__M5_1 vdd vdd vbp vbp bbp__M5
.ends

.subckt bbn__M2 a_50_n100# a_n50_n126# a_n108_n100# VSUBS
X0 a_50_n100# a_n50_n126# a_n108_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt bbn__M3 a_50_n100# a_n50_n126# a_n108_n100# VSUBS
X0 a_50_n100# a_n50_n126# a_n108_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt bbn__M1 a_50_n100# a_n50_n126# a_n108_n100# VSUBS
X0 a_50_n100# a_n50_n126# a_n108_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt bb__nmirr vres vbp vbn ibn vss
Xbbn__M2_30 vbp vbn vres vss bbn__M2
Xbbn__M3_0 ibn vbn vss vss bbn__M3
Xbbn__M2_31 vbp vbn vres vss bbn__M2
Xbbn__M2_20 vbp vbn vres vss bbn__M2
Xbbn__M3_1 ibn vbn vss vss bbn__M3
Xbbn__M2_21 vbp vbn vres vss bbn__M2
Xbbn__M2_10 vbp vbn vres vss bbn__M2
Xbbn__M2_22 vbp vbn vres vss bbn__M2
Xbbn__M2_11 vbp vbn vres vss bbn__M2
Xbbn__M2_23 vbp vbn vres vss bbn__M2
Xbbn__M2_12 vbp vbn vres vss bbn__M2
Xbbn__M1_0 vbn vbn vss vss bbn__M1
Xbbn__M1_1 vbn vbn vss vss bbn__M1
Xbbn__M2_13 vbp vbn vres vss bbn__M2
Xbbn__M2_24 vbp vbn vres vss bbn__M2
Xbbn__M1_2 vbn vbn vss vss bbn__M1
Xbbn__M2_14 vbp vbn vres vss bbn__M2
Xbbn__M2_25 vbp vbn vres vss bbn__M2
Xbbn__M1_3 vbn vbn vss vss bbn__M1
Xbbn__M2_26 vbp vbn vres vss bbn__M2
Xbbn__M2_15 vbp vbn vres vss bbn__M2
Xbbn__M1_4 vbn vbn vss vss bbn__M1
Xbbn__M2_16 vbp vbn vres vss bbn__M2
Xbbn__M2_27 vbp vbn vres vss bbn__M2
Xbbn__M1_5 vbn vbn vss vss bbn__M1
Xbbn__M2_28 vbp vbn vres vss bbn__M2
Xbbn__M2_17 vbp vbn vres vss bbn__M2
Xbbn__M1_6 vbn vbn vss vss bbn__M1
Xbbn__M2_29 vbp vbn vres vss bbn__M2
Xbbn__M2_18 vbp vbn vres vss bbn__M2
Xbbn__M1_7 vbn vbn vss vss bbn__M1
Xbbn__M2_19 vbp vbn vres vss bbn__M2
Xbbn__M2_0 vbp vbn vres vss bbn__M2
Xbbn__M2_1 vbp vbn vres vss bbn__M2
Xbbn__M2_2 vbp vbn vres vss bbn__M2
Xbbn__M2_3 vbp vbn vres vss bbn__M2
Xbbn__M2_4 vbp vbn vres vss bbn__M2
Xbbn__M2_5 vbp vbn vres vss bbn__M2
Xbbn__M2_6 vbp vbn vres vss bbn__M2
Xbbn__M2_7 vbp vbn vres vss bbn__M2
Xbbn__M2_8 vbp vbn vres vss bbn__M2
Xbbn__M2_9 vbp vbn vres vss bbn__M2
.ends

.subckt bb__r1 a_n194_n1132# a_n324_n1262# a_124_696# a_n194_696# a_124_n1132#
X0 a_124_696# a_124_n1132# a_n324_n1262# sky130_fd_pr__res_xhigh_po_0p35 l=7.12
X1 a_n194_696# a_n194_n1132# a_n324_n1262# sky130_fd_pr__res_xhigh_po_0p35 l=7.12
.ends

.subckt bb__M10 a_n100_n112# a_n158_n86# w_n194_n148# a_100_n86#
X0 a_100_n86# a_n100_n112# a_n158_n86# w_n194_n148# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
.ends

.subckt bb__M9 a_n100_n112# a_n158_n86# w_n194_n148# a_100_n86#
X0 a_100_n86# a_n100_n112# a_n158_n86# w_n194_n148# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
.ends

.subckt bb__M7 a_n33_91# a_30_n131# a_n88_n131#
X0 a_30_n131# a_n33_91# a_n88_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt bb__R2 a_124_n1282# a_124_846# a_n194_846# a_n194_n1282#
X0 a_124_846# a_124_n1282# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=8.62
X1 a_n194_846# a_n194_n1282# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=8.62
.ends

.subckt bb__M8 a_n33_91# a_30_n131# a_n88_n131#
X0 a_30_n131# a_n33_91# a_n88_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt bias_basis_current vsu ibp ibn vdd vss
Xbb__pmirr_0 bb__pmirr_0/vbn bb__pmirr_0/vbp ibp vdd bb__pmirr
Xbb__nmirr_0 bb__nmirr_0/vres bb__pmirr_0/vbp bb__pmirr_0/vbn ibn vss bb__nmirr
Xbb__r1_0 m1_1749_871# vss vss bb__nmirr_0/vres m1_1749_871# bb__r1
Xbb__M10_0 m2_490_5152# m2_97_3643# vdd m2_490_5152# bb__M10
Xbb__M9_0 vsu m2_490_5152# vdd vsu bb__M9
Xbb__M7_0 vsu vsu vss bb__M7
Xbb__R2_0 m2_97_3643# m1_322_845# m1_322_845# vdd bb__R2
Xbb__M8_0 vsu vdd bb__pmirr_0/vbn bb__M8
.ends

.subckt bg__cap c1_n1050_n1000# m3_n1150_n1100#
X0 c1_n1050_n1000# m3_n1150_n1100# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt bg__res a_n1613_1296# a_n455_n1732# a_n3157_n1732# a_1089_n1732# a_n1227_n1732#
+ a_317_1296# a_n2771_n1732# a_703_1296# a_2247_n1732# a_2247_1296# a_2633_1296# a_n69_n1732#
+ a_n3929_n1732# a_3791_n1732# a_n2385_1296# a_1861_n1732# a_703_n1732# a_n2771_1296#
+ a_n3929_1296# a_3405_n1732# a_n69_1296# a_n455_1296# a_n841_1296# a_n2385_n1732#
+ a_n1999_1296# a_n1999_n1732# a_3019_1296# a_3405_1296# a_n841_n1732# a_n3543_n1732#
+ a_3791_1296# a_1475_n1732# a_317_n1732# a_n1613_n1732# a_n3157_1296# a_3019_n1732#
+ a_1089_1296# a_n3543_1296# a_1475_1296# a_2633_n1732# a_1861_1296# a_n4059_n1862#
+ a_n1227_1296#
X0 a_317_1296# a_317_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X1 a_n69_1296# a_n69_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X2 a_1861_1296# a_1861_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X3 a_703_1296# a_703_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X4 a_n1227_1296# a_n1227_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X5 a_n2385_1296# a_n2385_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X6 a_2247_1296# a_2247_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X7 a_n1999_1296# a_n1999_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X8 a_n1613_1296# a_n1613_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X9 a_n2771_1296# a_n2771_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X10 a_2633_1296# a_2633_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X11 a_3791_1296# a_3791_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X12 a_n3157_1296# a_n3157_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X13 a_3019_1296# a_3019_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X14 a_n3543_1296# a_n3543_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X15 a_3405_1296# a_3405_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X16 a_n455_1296# a_n455_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X17 a_1089_1296# a_1089_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X18 a_n841_1296# a_n841_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X19 a_n3929_1296# a_n3929_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X20 a_1475_1296# a_1475_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
.ends

.subckt bgt__MN a_n108_n231# a_n210_n343# a_50_n231# a_n50_n257#
X0 a_50_n231# a_n50_n257# a_n108_n231# a_n210_n343# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt bgt__res a_n1996_n712# a_n3056_n712# a_124_276# a_n936_276# a_1714_276# a_1714_n712#
+ a_n2526_276# a_654_276# a_n1466_n712# a_n1466_276# a_n4116_n712# a_n4246_n842# a_3304_276#
+ a_2244_276# a_1184_n712# a_n4116_276# a_2774_n712# a_1184_276# a_n3056_276# a_n1996_276#
+ a_3834_276# a_n2526_n712# a_2774_276# a_654_n712# a_3834_n712# a_2244_n712# a_n936_n712#
+ a_n3586_276# a_n3586_n712# a_n406_276# a_124_n712# a_n406_n712# a_3304_n712#
X0 a_n1466_276# a_n1466_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X1 a_3834_276# a_3834_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X2 a_1714_276# a_1714_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X3 a_n936_276# a_n936_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X4 a_n3056_276# a_n3056_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X5 a_3304_276# a_3304_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X6 a_n406_276# a_n406_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X7 a_2774_276# a_2774_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X8 a_2244_276# a_2244_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X9 a_1184_276# a_1184_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X10 a_654_276# a_654_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X11 a_124_276# a_124_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X12 a_n2526_276# a_n2526_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X13 a_n1996_276# a_n1996_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X14 a_n4116_276# a_n4116_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X15 a_n3586_276# a_n3586_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
.ends

.subckt bg__trim m2_4223_3828# m2_800_5948# m2_640_4888# m2_4223_648# bgt__res_0/a_3834_n712#
+ m2_1120_8068# m2_480_3828# m2_4223_2768# m2_320_2768# m1_4339_1060# m1_1336_1060#
+ m2_4223_5948# m2_4223_8068# m2_160_1708# m1_3744_8480# m2_4223_4888# m2_4223_1708#
+ m2_960_7008# m2_0_648# VSUBS m2_4223_7008#
Xbgt__MN_0 m1_4339_1060# VSUBS m1_3744_8480# m2_4223_8068# bgt__MN
Xbgt__MN_1 m1_4339_1060# VSUBS m1_3323_1060# m2_4223_648# bgt__MN
Xbgt__MN_2 m1_4339_1060# VSUBS m1_3323_2120# m2_4223_1708# bgt__MN
Xbgt__MN_3 m1_4339_1060# VSUBS m1_3323_3180# m2_4223_2768# bgt__MN
Xbgt__MN_5 m1_4339_1060# VSUBS m1_3323_5300# m2_4223_4888# bgt__MN
Xbgt__MN_4 m1_4339_1060# VSUBS m1_3323_4240# m2_4223_3828# bgt__MN
Xbgt__MN_6 m1_1336_1060# VSUBS m1_1849_8480# m2_1120_8068# bgt__MN
Xbgt__MN_7 m1_4339_1060# VSUBS m1_3323_6360# m2_4223_5948# bgt__MN
Xbgt__MN_8 m1_4339_1060# VSUBS m1_3323_7420# m2_4223_7008# bgt__MN
Xbgt__MN_9 m1_1336_1060# VSUBS m1_1849_1060# m2_0_648# bgt__MN
Xbgt__MN_10 m1_1336_1060# VSUBS m1_1849_2120# m2_160_1708# bgt__MN
Xbgt__MN_11 m1_1336_1060# VSUBS m1_1849_3180# m2_320_2768# bgt__MN
Xbgt__MN_12 m1_1336_1060# VSUBS m1_1849_4240# m2_480_3828# bgt__MN
Xbgt__MN_13 m1_1336_1060# VSUBS m1_1849_5300# m2_640_4888# bgt__MN
Xbgt__MN_14 m1_1336_1060# VSUBS m1_1849_6360# m2_800_5948# bgt__MN
Xbgt__MN_15 m1_1336_1060# VSUBS m1_1849_7420# m2_960_7008# bgt__MN
Xbgt__res_0 m1_3323_6360# m1_3323_7420# m1_1849_4240# m1_1849_5300# m1_1849_3180#
+ m1_3323_2120# m1_1849_7420# m1_1849_4240# m1_3323_5300# m1_1849_6360# m1_3744_8480#
+ VSUBS m1_1849_1060# m1_1849_2120# m1_3323_3180# m1_1849_8480# m1_3323_1060# m1_1849_3180#
+ m1_1849_7420# m1_1849_6360# m1_1849_1060# m1_3323_6360# m1_1849_2120# m1_3323_3180#
+ bgt__res_0/a_3834_n712# m1_3323_2120# m1_3323_5300# m1_1849_8480# m1_3323_7420#
+ m1_1849_5300# m1_3323_4240# m1_3323_4240# m1_3323_1060# bgt__res
.ends

.subckt bgs__M3_M4 a_n287_n131# a_29_n157# a_229_n131# a_n229_n157# a_n389_n243# a_n29_n131#
X0 a_n29_n131# a_n229_n157# a_n287_n131# a_n389_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_229_n131# a_29_n157# a_n29_n131# a_n389_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt bgs__M5_M6 w_n425_n284# a_n287_n136# a_229_n136# a_29_n162# a_n29_n136# a_n229_n162#
X0 a_n29_n136# a_n229_n162# a_n287_n136# w_n425_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_229_n136# a_29_n162# a_n29_n136# w_n425_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt bgs__M7 a_100_n136# w_n296_n284# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n296_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bg__startup m2_545_805# VSUBS m1_453_173# bgs__M5_M6_0/w_n425_n284# m1_2508_588#
+ m2_1443_341# m1_1258_542# bgs__M7_0/w_n296_n284# bgs__M3_M4_0/a_n287_n131# bgs__M7_0/a_100_n136#
Xbgs__M3_M4_0 bgs__M3_M4_0/a_n287_n131# m2_545_805# m1_251_542# m1_251_542# VSUBS
+ m1_453_173# bgs__M3_M4
Xbgs__M5_M6_0 bgs__M5_M6_0/w_n425_n284# m1_251_542# m1_1258_542# m1_1258_542# m2_1443_341#
+ m1_1258_542# bgs__M5_M6
Xbgs__M7_0 bgs__M7_0/a_100_n136# bgs__M7_0/w_n296_n284# m1_1258_542# m1_2508_588#
+ bgs__M7
.ends

.subckt bg__M1_M2 a_n287_n436# a_n487_n462# w_n683_n584# a_229_n436# a_29_n462# a_n545_n436#
+ a_n29_n436# a_n229_n462# a_487_n436# a_287_n462#
X0 a_n287_n436# a_n487_n462# a_n545_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_487_n436# a_287_n462# a_229_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2 a_229_n436# a_29_n462# a_n29_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n29_n436# a_n229_n462# a_n287_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt bgpg__pnp a_26_26# w_153_153# a_330_330#
X0 a_26_26# w_153_153# a_330_330# sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544
.ends

.subckt bg__pnp_group eg eu VDD GND
Xbgpg__pnp_0 GND GND eg bgpg__pnp
Xbgpg__pnp_1 GND GND eg bgpg__pnp
Xbgpg__pnp_2 GND GND eg bgpg__pnp
Xbgpg__pnp_3 GND GND eg bgpg__pnp
Xbgpg__pnp_4 GND GND eg bgpg__pnp
Xbgpg__pnp_5 GND GND eg bgpg__pnp
Xbgpg__pnp_6 GND GND eu bgpg__pnp
Xbgpg__pnp_7 GND GND eg bgpg__pnp
Xbgpg__pnp_8 GND GND eg bgpg__pnp
.ends

.subckt bgfcpm__DUM w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcpm__M1 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcpm__MB2 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcpm__MB3 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfc__pmirr vbp1 diff vbn2 vdd
Xbgfcpm__DUM_3 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_28 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_17 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_4 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_0 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__DUM_29 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_18 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_5 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_1 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__DUM_19 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_6 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_2 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__DUM_7 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_3 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__M1_4 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__DUM_8 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_5 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__DUM_9 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_6 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__M1_7 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__M1_8 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__M1_9 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__MB2_0 vdd vdd vbp1 vbp1 bgfcpm__MB2
Xbgfcpm__M1_10 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__MB2_1 vdd vdd vbp1 vbp1 bgfcpm__MB2
Xbgfcpm__M1_11 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__MB2_2 vdd vbp1 vdd vbp1 bgfcpm__MB2
Xbgfcpm__M1_12 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__MB2_3 vdd vbp1 vdd vbp1 bgfcpm__MB2
Xbgfcpm__M1_13 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__M1_14 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__M1_15 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__DUM_30 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_20 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_31 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_21 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_10 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_22 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_11 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_0 vdd vbn2 vdd vbp1 bgfcpm__MB3
Xbgfcpm__DUM_23 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_12 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_1 vdd vdd vbn2 vbp1 bgfcpm__MB3
Xbgfcpm__DUM_24 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_13 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_2 vdd vbn2 vdd vbp1 bgfcpm__MB3
Xbgfcpm__DUM_0 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_25 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_14 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_3 vdd vdd vbn2 vbp1 bgfcpm__MB3
Xbgfcpm__DUM_1 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_15 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_26 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_2 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_16 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_27 vdd vdd vdd vdd bgfcpm__DUM
.ends

.subckt bgfcnm__M4 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcnm__M5 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcnm__MB5 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcnm__DUM a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfc__nmirr vbn1 out1n out1p vss
Xbgfcnm__M4_13 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_0 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_14 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_1 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_15 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_2 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_3 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_4 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_5 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_6 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_7 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_8 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M5_10 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__MB5_0 vbn1 vbn1 vss vss bgfcnm__MB5
Xbgfcnm__M4_9 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__MB5_1 vss vbn1 vbn1 vss bgfcnm__MB5
Xbgfcnm__M5_11 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__M5_12 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__MB5_2 vss vbn1 vbn1 vss bgfcnm__MB5
Xbgfcnm__DUM_40 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_13 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__MB5_3 vbn1 vbn1 vss vss bgfcnm__MB5
Xbgfcnm__DUM_41 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_30 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_42 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_31 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_14 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_20 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_15 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_21 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_32 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_43 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_0 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_10 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_33 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_22 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_11 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_1 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_23 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_34 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_12 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_2 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_0 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_35 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_24 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_13 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_3 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_1 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_36 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_25 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_14 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_4 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_2 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_37 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_26 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_15 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_5 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_3 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_38 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_27 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_16 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_6 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_4 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_39 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_28 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_17 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_7 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_5 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_29 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_18 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_8 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_6 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_9 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_19 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_7 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__M5_8 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__M5_9 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__M4_10 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_11 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_12 vss vbn1 out1n vss bgfcnm__M4
.ends

.subckt bgfccpt__DUM a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpt__M11 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpt__M10 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfc__casp_top vdd nd11 nd10 mirr m1_458_30#
Xbgfccpt__DUM_7 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_8 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__M11_0 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_9 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_1 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_20 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_2 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_21 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_10 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_3 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_22 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_11 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_4 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_12 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_23 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_5 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_13 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_6 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_14 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__M11_7 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_15 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_16 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_17 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_18 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_19 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__M10_0 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__M10_1 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_2 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_3 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_4 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__M10_5 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_6 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__M10_7 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__DUM_0 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__DUM_1 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_2 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_3 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_4 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_5 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_6 vdd vdd m1_458_30# vdd bgfccpt__DUM
.ends

.subckt bgfccnt__M6 a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfccnt__DUM a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfccnt__M7 a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfccnt__MB4 a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfc__casn_top vbn2 vbn1 out mirr out1n out1p VSUBS
Xbgfccnt__M6_0 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__M6_1 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__M6_2 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__M6_3 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__M6_4 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__DUM_0 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M6_5 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__DUM_1 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
Xbgfccnt__M6_6 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__DUM_2 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M6_7 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__DUM_3 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_4 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_5 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_6 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_7 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_8 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
Xbgfccnt__DUM_9 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M7_0 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__M7_1 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__M7_2 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__DUM_20 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_0 vbn1 vbn2 vbn2 VSUBS bgfccnt__MB4
Xbgfccnt__M7_3 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__DUM_10 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_21 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_1 vbn1 vbn2 vbn2 VSUBS bgfccnt__MB4
Xbgfccnt__M7_4 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__DUM_11 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_22 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_2 vbn2 vbn2 vbn1 VSUBS bgfccnt__MB4
Xbgfccnt__M7_5 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__DUM_12 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_23 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_3 vbn2 vbn2 vbn1 VSUBS bgfccnt__MB4
Xbgfccnt__M7_6 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__DUM_13 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_24 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M7_7 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__DUM_14 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_25 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_26 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_15 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
Xbgfccnt__DUM_16 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_27 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_17 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_18 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_19 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
.ends

.subckt bgfcdpp__M3 w_n194_n498# a_100_n436# a_n158_n436# a_n100_n462#
X0 a_100_n436# a_n100_n462# a_n158_n436# w_n194_n498# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt bgfcdpp__M2 w_n194_n498# a_100_n436# a_n158_n436# a_n100_n462#
X0 a_100_n436# a_n100_n462# a_n158_n436# w_n194_n498# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt bgfcdpp__DUM w_n194_n498# a_100_n436# a_n158_n436# a_n100_n462#
X0 a_100_n436# a_n100_n462# a_n158_n436# w_n194_n498# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt bgfc__diffpair_p inp inn diff out1p out1n vdd
Xbgfcdpp__M3_0 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_1 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M3_2 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_3 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M3_4 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_5 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M3_6 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_7 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M2_0 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__M2_1 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_2 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__M2_3 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_4 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__M2_5 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_6 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_7 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__DUM_0 vdd diff diff diff bgfcdpp__DUM
Xbgfcdpp__DUM_1 vdd diff diff diff bgfcdpp__DUM
Xbgfcdpp__DUM_2 vdd diff diff diff bgfcdpp__DUM
Xbgfcdpp__DUM_3 vdd diff diff diff bgfcdpp__DUM
.ends

.subckt bgfccpb__M8 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpb__M9 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpb__DUM a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpb__MB1 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfc__casp_bot out nd11 nd10 mirr bias vbp1 m1_458_17#
Xbgfccpb__M8_0 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M8_1 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_2 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M8_3 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_4 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_5 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M8_6 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_7 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M9_0 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__M9_1 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__DUM_0 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__M9_2 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__MB1_0 vbp1 bias m1_458_17# bias bgfccpb__MB1
Xbgfccpb__M9_3 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__DUM_1 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__MB1_1 vbp1 bias m1_458_17# bias bgfccpb__MB1
Xbgfccpb__DUM_2 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__M9_4 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__MB1_2 bias bias m1_458_17# vbp1 bgfccpb__MB1
Xbgfccpb__M9_5 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__DUM_3 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_20 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__MB1_3 bias bias m1_458_17# vbp1 bgfccpb__MB1
Xbgfccpb__DUM_4 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__M9_6 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__DUM_21 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_10 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__M9_7 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__DUM_5 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_22 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_11 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_6 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_23 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_12 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__DUM_7 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_24 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_13 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_8 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_14 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_25 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__DUM_9 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_26 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_15 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_16 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__DUM_27 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_17 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_18 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_19 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
.ends

.subckt bg__se_folded_cascode_p vbn1 vbp1 diff out1p out1n mirr vbn2 nd10 nd11 out
+ vdd bias vsub inp inn vss
Xbgfc__pmirr_0 vbp1 diff vbn2 vdd bgfc__pmirr
Xbgfc__nmirr_0 vbn1 out1n out1p vss bgfc__nmirr
Xbgfc__casp_top_0 vdd nd11 nd10 mirr vdd bgfc__casp_top
Xbgfc__casn_top_0 vbn2 vbn1 out mirr out1n out1p vss bgfc__casn_top
Xbgfc__diffpair_p_0 inp inn diff out1p out1n vdd bgfc__diffpair_p
Xbgfc__casp_bot_0 out nd11 nd10 mirr bias vbp1 vdd bgfc__casp_bot
.ends

.subckt bandgap_cw vbg trim[15] trim[13] trim[11] trim[9] trim[7] trim[5] trim[3]
+ trim[1] trim[0] trim[2] trim[4] trim[6] trim[8] trim[10] trim[12] trim[14] bias
+ vdd vsub vss
Xbg__cap_3 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_4 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__res_0 m1_32787_8825# m1_32015_12378# m1_35489_12378# m1_30085_12378# m1_33559_12378#
+ m1_30857_8825# m1_35103_12378# m1_31243_9043# m1_30085_12378# m1_29699_9043# m1_29699_9043#
+ m2_32390_12378# m1_35103_12378# m1_28541_12378# m1_34717_9043# m1_30471_12378# m1_31629_12378#
+ m1_34717_9043# m1_33977_7455# m1_28927_12378# bg__se_folded_cascode_p_0/inp m1_32787_8825#
+ m1_33173_9043# m1_33559_12378# m1_34331_8825# m1_33945_12378# m1_29313_8825# bg__se_folded_cascode_p_0/inp
+ m1_31629_12378# m1_35489_12378# bg__pnp_group_0/eu m1_30471_12378# m1_32015_12378#
+ m1_33945_12378# m1_34331_8825# m1_28927_12378# m1_31243_9043# vbg m1_30857_8825#
+ m1_28541_12378# m1_29313_8825# vss m1_33173_9043# bg__res
Xbg__cap_5 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_6 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_7 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_8 vdd vss bg__cap
Xbg__trim_0 trim[7] trim[10] trim[8] trim[1] bg__pnp_group_0/eg trim[14] trim[6] trim[5]
+ trim[4] bg__pnp_group_0/eg bg__pnp_group_0/eg trim[11] trim[15] trim[2] m2_32390_12378#
+ trim[9] trim[3] trim[12] trim[0] vss trim[13] bg__trim
Xbg__cap_9 vdd vss bg__cap
Xbg__startup_0 vbg vss vss vdd vdd vdd vdd vdd bg__se_folded_cascode_p_0/out vss bg__startup
Xbg__M1_M2_0 vbg bg__se_folded_cascode_p_0/out vdd m1_33977_7455# bg__se_folded_cascode_p_0/out
+ vdd vdd bg__se_folded_cascode_p_0/out vdd bg__se_folded_cascode_p_0/out bg__M1_M2
Xbg__pnp_group_0 bg__pnp_group_0/eg bg__pnp_group_0/eu vdd vss bg__pnp_group
Xbg__cap_10 vdd vss bg__cap
Xbg__se_folded_cascode_p_0 bg__se_folded_cascode_p_0/vbn1 bg__se_folded_cascode_p_0/vbp1
+ bg__se_folded_cascode_p_0/diff bg__se_folded_cascode_p_0/out1p bg__se_folded_cascode_p_0/out1n
+ bg__se_folded_cascode_p_0/mirr bg__se_folded_cascode_p_0/vbn2 bg__se_folded_cascode_p_0/nd10
+ bg__se_folded_cascode_p_0/nd11 bg__se_folded_cascode_p_0/out vdd bias vsub bg__se_folded_cascode_p_0/inp
+ bg__pnp_group_0/eu vss bg__se_folded_cascode_p
Xbg__cap_0 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_1 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_2 bg__se_folded_cascode_p_0/out vss bg__cap
.ends

.subckt sky130_cw_ip__bandgap trim[0] trim[4] trim[6] trim[10] trim[12] trim[14] trim[15]
+ trim[13] trim[11] trim[7] trim[5] trim[3] trim[1] trim[2] vbg trim[8] trim[9] vdd
+ vsub vss
Xbias_basis_current_0 bias_basis_current_0/vsu bias_basis_current_0/ibp bandgap_cw_0/bias
+ vdd vss bias_basis_current
Xbandgap_cw_0 vbg trim[15] trim[13] trim[11] trim[9] trim[7] trim[5] trim[3] trim[1]
+ trim[0] trim[2] trim[4] trim[6] trim[8] trim[10] trim[12] trim[14] bandgap_cw_0/bias
+ vdd vsub vss bandgap_cw
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RBNV2H a_n287_n188# a_n29_n100# a_345_n188# a_n445_n188#
+ a_n187_n100# a_503_n188# a_n603_n188# a_n345_n100# a_129_n100# a_n503_n100# a_n661_n100#
+ a_287_n100# a_445_n100# a_29_n188# a_n129_n188# a_603_n100# a_187_n188# a_n795_n322#
X0 a_445_n100# a_345_n188# a_287_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_603_n100# a_503_n188# a_445_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X2 a_129_n100# a_29_n188# a_n29_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n187_n100# a_n287_n188# a_n345_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n345_n100# a_n445_n188# a_n503_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n503_n100# a_n603_n188# a_n661_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X6 a_n29_n100# a_n129_n188# a_n187_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_287_n100# a_187_n188# a_129_n100# a_n795_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_ZB8LT7 a_1560_11084# a_48_n11516# a_n1972_n11646#
+ a_804_n11516# a_1560_n11516# a_48_11084# a_n330_11084# a_n708_11084# a_426_n11516#
+ a_n1086_11084# a_n1464_11084# a_1182_n11516# a_n1842_11084# a_n330_n11516# a_n1842_n11516#
+ a_n708_n11516# a_426_11084# a_804_11084# a_n1464_n11516# a_1182_11084# a_n1086_n11516#
X0 a_804_11084# a_804_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X1 a_n1464_11084# a_n1464_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X2 a_426_11084# a_426_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X3 a_n708_11084# a_n708_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X4 a_1560_11084# a_1560_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X5 a_n1086_11084# a_n1086_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X6 a_n1842_11084# a_n1842_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X7 a_n330_11084# a_n330_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X8 a_1182_11084# a_1182_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
X9 a_48_11084# a_48_n11516# a_n1972_n11646# sky130_fd_pr__res_xhigh_po_1p41 l=111
.ends

.subckt rc_osc_por dvdd out ena dvss
Xsky130_fd_pr__pfet_01v8_MA8JJJ_0 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_MA8JJJ
Xsky130_fd_pr__res_xhigh_po_1p41_ZB8LT7_0 m1_25146_n1894# m1_2270_n760# dvss m1_2270_n1516#
+ in m1_25146_n382# m1_25146_n382# m1_25146_374# m1_2270_n760# m1_25146_374# m1_25146_1130#
+ m1_2270_n1516# m1_25146_1130# m1_2270_n4# vr m1_2270_n4# m1_25146_n1138# m1_25146_n1138#
+ m1_2270_752# m1_25146_n1894# m1_2270_752# sky130_fd_pr__res_xhigh_po_1p41_ZB8LT7
Xsky130_fd_pr__pfet_01v8_LAUYMQ_0 dvdd dvdd vr ena_b out dvdd sky130_fd_pr__pfet_01v8_LAUYMQ
Xsky130_fd_pr__pfet_01v8_C64SS5_0 m dvdd dvdd dvdd in in in m in dvdd in m dvdd in
+ sky130_fd_pr__pfet_01v8_C64SS5
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 in dvdd dvdd ena sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_C68ZY6_0 out n n dvdd dvdd m n n out m n dvdd dvdd dvdd m
+ m sky130_fd_pr__pfet_01v8_C68ZY6
Xsky130_fd_pr__pfet_01v8_C6GQGA_0 dvdd dvdd ena_b ena sky130_fd_pr__pfet_01v8_C6GQGA
Xsky130_fd_pr__pfet_01v8_9QCJ55_0 m m n n n dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_9QCJ55
Xsky130_fd_pr__pfet_01v8_MLERZ7_0 vr ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_MLERZ7
X0 dvss dvss m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 m n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 dvss ena ena_b dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 out ena vr dvss sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X4 dvss dvss n dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 dvss in m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 n m dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 dvss dvss out dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X8 m in dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X9 vr dvss dvss dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X10 out n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X3 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X8 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X11 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X15 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X16 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X18 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X19 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X20 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X21 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X22 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X23 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X24 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X25 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X26 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X27 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X28 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X29 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X30 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X31 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt por_ana otrip_decoded[7] otrip_decoded[5] otrip_decoded[3] otrip_decoded[1]
+ vbg_1v2 itest ibg_200n dvdd dcomp isrc_sel pwup_filt osc_ck osc_ena porb_h por porb
+ comparator_1/vt force_pdnb otrip_decoded[4] comparator_0/vt otrip_decoded[2] por_unbuf
+ avdd vin otrip_decoded[6] otrip_decoded[0] avss dvss
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_4_4/Y dvss dvss dvdd dvdd por sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hvl__lsbufhv2lv_1_0 dcomp3v3 dvdd dvss dvss avdd avdd vl sky130_fd_sc_hvl__lsbufhv2lv_1
Xsky130_fd_sc_hvl__lsbufhv2lv_1_1 dcomp3v3uv dvdd dvss dvss avdd avdd sky130_fd_sc_hvl__lsbufhv2lv_1_1/X
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xrstring_mux_0 vin ibias_gen_0/ena rstring_mux_0/otrip_decoded_avdd[7] rstring_mux_0/otrip_decoded_avdd[6]
+ rstring_mux_0/otrip_decoded_avdd[5] rstring_mux_0/otrip_decoded_avdd[4] rstring_mux_0/otrip_decoded_avdd[3]
+ rstring_mux_0/otrip_decoded_avdd[2] rstring_mux_0/otrip_decoded_avdd[1] rstring_mux_0/vtrip_decoded_avdd[7]
+ rstring_mux_0/vtrip_decoded_avdd[6] rstring_mux_0/vtrip_decoded_avdd[5] rstring_mux_0/vtrip_decoded_avdd[4]
+ rstring_mux_0/vtrip_decoded_avdd[3] rstring_mux_0/vtrip_decoded_avdd[2] rstring_mux_0/vtrip_decoded_avdd[1]
+ rstring_mux_0/vtrip_decoded_avdd[0] comparator_0/vinn rstring_mux_0/vtop rstring_mux_0/otrip_decoded_avdd[0]
+ avdd avss rstring_mux
Xsky130_fd_sc_hvl__inv_4_0 sky130_fd_sc_hvl__inv_4_0/A avss avss avdd avdd sky130_fd_sc_hvl__inv_4_0/Y
+ sky130_fd_sc_hvl__inv_4
Xsky130_fd_sc_hd__inv_4_0 schmitt_trigger_0/out dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_0/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_1 sky130_fd_sc_hd__inv_4_2/Y dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_2 por_unbuf dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_2/Y
+ sky130_fd_sc_hd__inv_4
Xschmitt_trigger_0 schmitt_trigger_0/in schmitt_trigger_0/out dvdd dvss schmitt_trigger
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] otrip_decoded[0] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] otrip_decoded[1] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] otrip_decoded[2] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] otrip_decoded[3] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2] otrip_decoded[4] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2] otrip_decoded[5] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3] otrip_decoded[6] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3] otrip_decoded[7] dvdd dvss dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[0]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[1]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[2]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[3]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[4]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[5]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[6]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7] dvss dvdd dvss dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[7]
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8] force_pdnb dvdd dvss dvss avdd avdd ibias_gen_0/ena
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8] isrc_sel dvdd dvss dvss avdd avdd ibias_gen_0/isrc_sel
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hd__inv_4_3 vl dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hvl__lsbuflv2hv_1_1 por_unbuf dvdd dvss dvss avdd avdd sky130_fd_sc_hvl__inv_1_0/A
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hd__inv_4_4 por_unbuf dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_4/Y
+ sky130_fd_sc_hd__inv_4
Xrc_osc_por_0 dvdd osc_ck osc_ena dvss rc_osc_por
Xsky130_fd_sc_hvl__inv_16_0 sky130_fd_sc_hvl__inv_4_0/Y avss avss avdd avdd porb_h
+ sky130_fd_sc_hvl__inv_16
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_n11325_2001# m1_n11325_2001# m1_n12081_2001#
+ m1_n10191_9400# m1_n13971_9400# m1_n14349_2001# m1_n12081_2001# vl m1_n12837_2001#
+ m1_n8301_2001# m1_n12837_2001# avss m1_n9435_9400# m1_n10947_9400# m1_n13215_9400#
+ m1_n13215_9400# m1_n8679_9400# m1_n10569_2001# m1_n9435_9400# m1_n13971_9400# m1_n10569_2001#
+ m1_n14727_9400# m1_n8301_2001# m1_n10947_9400# m1_n13593_2001# schmitt_trigger_0/in
+ m1_n11703_9400# m1_n8679_9400# m1_n9813_2001# m1_n9057_2001# m1_n9813_2001# m1_n7923_9400#
+ m1_n12459_9400# m1_n11703_9400# m1_n13593_2001# m1_n14727_9400# m1_n10191_9400#
+ m1_n14349_2001# m1_n9057_2001# m1_n7923_9400# m1_n12459_9400# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 schmitt_trigger_0/in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xibias_gen_0 ibias_gen_0/ibias0 itest ibias_gen_0/ibias1 ibg_200n vbg_1v2 ibias_gen_0/isrc_sel
+ ibias_gen_0/ena ibias_gen_0/ve avss avdd ibias_gen
Xsky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 avss avss ibias_gen_0/ve sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 m=1
Xsky130_fd_sc_hvl__inv_1_0 sky130_fd_sc_hvl__inv_1_0/A avss avss avdd avdd sky130_fd_sc_hvl__inv_4_0/A
+ sky130_fd_sc_hvl__inv_1
Xcomparator_0 ibias_gen_0/ibias1 dcomp3v3uv avss comparator_0/vinn vbg_1v2 avss comparator_0/vt
+ avdd comparator
Xcomparator_1 ibias_gen_0/ibias0 dcomp3v3 ibias_gen_0/ena vbg_1v2 vin avss comparator_1/vt
+ avdd comparator
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_4_0/Y dvss dvss dvdd dvdd pwup_filt
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_4_1/Y dvss dvss dvdd dvdd porb sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_4_3/Y dvss dvss dvdd dvdd dcomp sky130_fd_sc_hd__inv_16
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05985 ps=0.705 w=0.42 l=0.15
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt por_dig force_dis_rc_osc force_short_oneshot osc_ck osc_ena otrip[0] otrip[1]
+ otrip[2] otrip_decoded[0] otrip_decoded[1] otrip_decoded[2] otrip_decoded[3] otrip_decoded[4]
+ otrip_decoded[5] otrip_decoded[6] otrip_decoded[7] por_timed_out por_unbuf pwup_filt
+ startup_timed_out force_pdn force_pdnb force_ena_rc_osc VPWR VGND
XFILLER_0_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_131_ clknet_1_0__leaf_osc_ck net29 net8 VGND VGND VPWR VPWR cnt_rsb sky130_fd_sc_hd__dfrtp_1
X_062_ net7 net6 net5 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__nor3b_1
X_114_ clknet_1_0__leaf_osc_ck net36 net24 VGND VGND VPWR VPWR cnt_st\[1\] sky130_fd_sc_hd__dfrtp_1
Xoutput20 net20 VGND VGND VPWR VPWR por_unbuf sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ clknet_1_0__leaf_osc_ck net27 net8 VGND VGND VPWR VPWR cnt_rsb_stg1 sky130_fd_sc_hd__dfrtp_1
X_113_ clknet_1_0__leaf_osc_ck _000_ net24 VGND VGND VPWR VPWR cnt_st\[0\] sky130_fd_sc_hd__dfrtp_1
X_061_ net7 net6 net5 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__nor3_1
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput21 net23 VGND VGND VPWR VPWR startup_timed_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
X_060_ net22 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__inv_2
Xhold10 cnt_por\[5\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
X_112_ net31 _026_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput11 net11 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR force_pdnb sky130_fd_sc_hd__buf_2
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_111_ _026_ _027_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold11 cnt_por\[1\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ cnt_por\[8\] net23 net22 _024_ net42 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a41o_1
Xhold12 cnt_por\[7\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput13 net13 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_0_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold13 cnt_por\[2\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_099_ _034_ _049_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__and2_1
Xhold14 cnt_st\[2\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
XFILLER_0_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ cnt_por\[4\] _049_ cnt_por\[5\] VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21oi_1
Xhold15 cnt_por\[9\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
X_097_ net26 _036_ _018_ _017_ net34 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o32a_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ cnt_por\[4\] _049_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ cnt_st\[3\] net26 _039_ _040_ _030_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__o311a_1
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_095_ net33 _048_ _017_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o21ba_1
Xoutput19 net19 VGND VGND VPWR VPWR por_timed_out sky130_fd_sc_hd__buf_2
X_078_ net26 _039_ cnt_st\[3\] VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_094_ net4 _049_ _035_ net21 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o211a_1
X_129_ clknet_1_0__leaf_osc_ck _016_ net24 VGND VGND VPWR VPWR cnt_por\[10\] sky130_fd_sc_hd__dfrtp_1
X_077_ _038_ _039_ net26 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ cnt_por\[1\] cnt_por\[0\] cnt_por\[3\] cnt_por\[2\] VGND VGND VPWR VPWR _049_
+ sky130_fd_sc_hd__and4_1
Xfanout22 _035_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_076_ cnt_st\[0\] cnt_st\[1\] cnt_st\[2\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__and3_1
Xinput1 force_dis_rc_osc VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_128_ clknet_1_0__leaf_osc_ck _015_ net24 VGND VGND VPWR VPWR cnt_por\[9\] sky130_fd_sc_hd__dfrtp_1
X_059_ _031_ _032_ _033_ _034_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or4bb_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout23 net21 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xinput2 force_ena_rc_osc VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_092_ cnt_por\[2\] net21 net22 _045_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and4_1
X_058_ cnt_por\[5\] cnt_por\[4\] VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__and2_1
X_127_ clknet_1_0__leaf_osc_ck _014_ net24 VGND VGND VPWR VPWR cnt_por\[8\] sky130_fd_sc_hd__dfrtp_1
X_075_ cnt_st\[0\] cnt_st\[1\] net41 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a21oi_1
Xfanout24 net28 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
X_091_ _043_ _046_ _047_ _036_ net40 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a32o_1
X_074_ cnt_st\[0\] net35 net23 _037_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a211oi_1
Xinput3 force_pdn VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_057_ cnt_por\[9\] cnt_por\[8\] VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__and2_1
X_126_ clknet_1_0__leaf_osc_ck _013_ net24 VGND VGND VPWR VPWR cnt_por\[7\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_109_ net23 _033_ net22 _024_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and4_1
Xfanout25 net28 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
X_090_ cnt_por\[2\] _045_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nand2_1
Xinput4 force_short_oneshot VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_0_5_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_125_ clknet_1_0__leaf_osc_ck _012_ net24 VGND VGND VPWR VPWR cnt_por\[6\] sky130_fd_sc_hd__dfrtp_1
X_073_ cnt_st\[0\] cnt_st\[1\] net26 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__o21bai_1
X_056_ cnt_por\[0\] cnt_por\[3\] cnt_por\[2\] cnt_por\[1\] VGND VGND VPWR VPWR _032_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_130__27 VGND VGND VPWR VPWR net27 _130__27/LO sky130_fd_sc_hd__conb_1
X_108_ net32 _025_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__xor2_1
Xfanout26 net4 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 otrip[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_072_ net26 net23 cnt_st\[0\] VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__or3b_1
X_124_ clknet_1_0__leaf_osc_ck _011_ net24 VGND VGND VPWR VPWR cnt_por\[5\] sky130_fd_sc_hd__dfrtp_1
X_055_ cnt_por\[7\] cnt_por\[6\] cnt_por\[10\] VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_6_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_107_ net39 _023_ _025_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__o21ba_1
X_071_ _036_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 otrip[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_55 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_054_ net23 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
X_123_ clknet_1_0__leaf_osc_ck _010_ net24 VGND VGND VPWR VPWR cnt_por\[4\] sky130_fd_sc_hd__dfrtp_1
X_106_ net23 net22 _024_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_070_ net23 net22 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 otrip[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_122_ clknet_1_1__leaf_osc_ck _009_ net25 VGND VGND VPWR VPWR cnt_por\[3\] sky130_fd_sc_hd__dfrtp_1
X_053_ cnt_st\[1\] _029_ cnt_st\[0\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and3b_1
XFILLER_0_2_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_105_ cnt_por\[7\] cnt_por\[6\] _034_ _049_ net26 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a41o_1
XFILLER_0_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
Xinput8 pwup_filt VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_121_ clknet_1_1__leaf_osc_ck _008_ net25 VGND VGND VPWR VPWR cnt_por\[2\] sky130_fd_sc_hd__dfrtp_1
X_104_ cnt_por\[6\] net23 net22 _020_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__and4_1
X_052_ cnt_st\[3\] cnt_st\[4\] cnt_st\[5\] cnt_st\[2\] VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ clknet_1_1__leaf_osc_ck _007_ net25 VGND VGND VPWR VPWR cnt_por\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_051_ net1 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
X_103_ cnt_por\[6\] _036_ _043_ _022_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_13_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 cnt_rsb VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
X_102_ cnt_por\[6\] _020_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__xor2_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
X_050_ net3 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__inv_2
Xhold2 cnt_rsb_stg1 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_101_ _043_ _021_ net37 net20 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 cnt_st\[5\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
X_100_ _019_ _020_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold4 cnt_por\[10\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold5 cnt_por\[8\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_089_ cnt_por\[2\] _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__or2_1
Xhold6 cnt_por\[3\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ _043_ _045_ _044_ net38 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__o2bb2a_1
Xhold7 cnt_por\[4\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ cnt_por\[1\] cnt_por\[0\] VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__and2_1
Xhold8 cnt_st\[1\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
X_086_ cnt_por\[0\] net26 net21 net22 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__o211a_1
Xhold9 _001_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
X_069_ net8 _028_ net22 net2 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__a31o_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _043_ _036_ cnt_por\[0\] VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__mux2_1
X_068_ net7 net6 net5 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__and3_1
X_084_ net26 net23 net22 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_067_ net5 net6 net7 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3b_1
X_119_ clknet_1_1__leaf_osc_ck _006_ net24 VGND VGND VPWR VPWR cnt_por\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_083_ net30 _041_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__xor2_1
X_118_ clknet_1_1__leaf_osc_ck _005_ net25 VGND VGND VPWR VPWR cnt_st\[5\] sky130_fd_sc_hd__dfrtp_1
X_066_ net6 net5 net7 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_16_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_082_ _041_ _042_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nor2_1
X_065_ net6 net5 net7 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_4_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_117_ clknet_1_1__leaf_osc_ck _004_ net25 VGND VGND VPWR VPWR cnt_st\[4\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_081_ cnt_st\[4\] _040_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_064_ net7 net6 net5 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__and3b_1
X_116_ clknet_1_1__leaf_osc_ck _003_ net25 VGND VGND VPWR VPWR cnt_st\[3\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_080_ net26 _039_ cnt_st\[3\] cnt_st\[4\] VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ net7 net5 net6 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor3b_1
X_115_ clknet_1_0__leaf_osc_ck _002_ net25 VGND VGND VPWR VPWR cnt_st\[2\] sky130_fd_sc_hd__dfrtp_1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_X6E435 a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MUZ6AA a_n287_n188# a_761_n100# a_n29_n100# a_345_n188#
+ a_n953_n322# a_n445_n188# a_n187_n100# a_503_n188# a_n819_n100# a_n603_n188# a_n345_n100#
+ a_661_n188# a_n761_n188# a_129_n100# a_n503_n100# a_n661_n100# a_287_n100# a_445_n100#
+ a_29_n188# a_n129_n188# a_603_n100# a_187_n188#
X0 a_445_n100# a_345_n188# a_287_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_603_n100# a_503_n188# a_445_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n661_n100# a_n761_n188# a_n819_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_129_n100# a_29_n188# a_n29_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n187_n100# a_n287_n188# a_n345_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n345_n100# a_n445_n188# a_n503_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n503_n100# a_n603_n188# a_n661_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n29_n100# a_n129_n188# a_n187_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_761_n100# a_661_n188# a_603_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X9 a_287_n100# a_187_n188# a_129_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_ajc_ip__por avdd dvdd vbg_1v2 otrip[2] otrip[1] otrip[0] force_pdn
+ force_ena_rc_osc force_short_oneshot isrc_sel ibg_200n vin porb_h porb por osc_ck
+ pwup_filt itest startup_timed_out por_timed_out force_dis_rc_osc dcomp por_ana_0/comparator_1/vt
+ por_ana_0/comparator_0/vt avss dvss
Xsky130_fd_pr__nfet_g5v0d10v5_RBNV2H_0 dvss dvss dvss dvss force_ena_rc_osc dvss dvss
+ dvss force_dis_rc_osc vbg_1v2 dvss dvss force_pdn dvss dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_RBNV2H
Xpor_ana_0 por_dig_0/otrip_decoded[7] por_dig_0/otrip_decoded[5] por_dig_0/otrip_decoded[3]
+ por_dig_0/otrip_decoded[1] vbg_1v2 itest ibg_200n dvdd dcomp isrc_sel pwup_filt
+ osc_ck por_dig_0/osc_ena porb_h por porb por_ana_0/comparator_1/vt por_dig_0/force_pdnb
+ por_dig_0/otrip_decoded[4] por_ana_0/comparator_0/vt por_dig_0/otrip_decoded[2]
+ por_dig_0/por_unbuf avdd vin por_dig_0/otrip_decoded[6] por_dig_0/otrip_decoded[0]
+ avss dvss por_ana
Xpor_dig_0 force_dis_rc_osc force_short_oneshot osc_ck por_dig_0/osc_ena otrip[0]
+ otrip[1] otrip[2] por_dig_0/otrip_decoded[0] por_dig_0/otrip_decoded[1] por_dig_0/otrip_decoded[2]
+ por_dig_0/otrip_decoded[3] por_dig_0/otrip_decoded[4] por_dig_0/otrip_decoded[5]
+ por_dig_0/otrip_decoded[6] por_dig_0/otrip_decoded[7] por_timed_out por_dig_0/por_unbuf
+ pwup_filt startup_timed_out force_pdn por_dig_0/force_pdnb force_ena_rc_osc dvdd
+ dvss por_dig
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_0 dvss vin dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_pr__nfet_g5v0d10v5_MUZ6AA_0 dvss dvss otrip[2] dvss dvss dvss dvss dvss
+ dvss dvss otrip[1] dvss dvss dvss dvss otrip[0] force_short_oneshot dvss dvss dvss
+ isrc_sel dvss sky130_fd_pr__nfet_g5v0d10v5_MUZ6AA
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_4V4BDM a_n29_n50# a_n187_n50# w_n387_n347# a_29_n147#
+ a_n129_n147# a_129_n50#
X0 a_129_n50# a_29_n147# a_n29_n50# w_n387_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_n50# a_n129_n147# a_n187_n50# w_n387_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8T5BGA a_n187_n136# a_129_n136# w_n387_n362#
+ a_29_n162# a_n129_n162# a_n29_n136#
X0 a_n29_n136# a_n129_n162# a_n187_n136# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_129_n136# a_29_n162# a_n29_n136# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_C5EREZ a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_S48KL6 a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt level_shifter_up VDD_HV x_lv x_hv xb_hv VDD_LV VSUBS m1_380_440# GND_HV
Xsky130_fd_pr__pfet_g5v0d10v5_4V4BDM_0 VDD_HV xb_hv VDD_HV xb_hv x_hv x_hv sky130_fd_pr__pfet_g5v0d10v5_4V4BDM
Xsky130_fd_pr__pfet_g5v0d10v5_8T5BGA_0 m1_380_440# m1_380_440# VDD_LV x_lv x_lv VDD_LV
+ sky130_fd_pr__pfet_g5v0d10v5_8T5BGA
Xsky130_fd_pr__nfet_g5v0d10v5_C5EREZ_0 m1_380_440# VSUBS VSUBS x_lv sky130_fd_pr__nfet_g5v0d10v5_C5EREZ
Xsky130_fd_pr__nfet_g5v0d10v5_S48KL6_0 GND_HV GND_HV x_hv xb_hv x_lv m1_380_440# sky130_fd_pr__nfet_g5v0d10v5_S48KL6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RUG6CB a_n400_n497# a_400_n400# w_n658_n697#
+ a_n458_n400#
X0 a_400_n400# a_n400_n497# a_n458_n400# w_n658_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_M7X63G a_150_n800# a_n208_n800# a_n150_n888#
+ a_n342_n1022#
X0 a_150_n800# a_n150_n888# a_n208_n800# a_n342_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_REE66T a_n487_n497# a_487_n400# a_n29_n400# a_545_n497#
+ a_n803_n400# a_29_n497# a_n287_n400# a_n1061_n400# a_n745_n497# a_803_n497# a_745_n400#
+ a_n229_n497# a_287_n497# a_n1003_n497# a_229_n400# a_n545_n400# w_n1261_n697# a_1003_n400#
X0 a_n545_n400# a_n745_n497# a_n803_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_n803_n400# a_n1003_n497# a_n1061_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2 a_n287_n400# a_n487_n497# a_n545_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_1003_n400# a_803_n497# a_745_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X4 a_487_n400# a_287_n497# a_229_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_745_n400# a_545_n497# a_487_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n29_n400# a_n229_n497# a_n287_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_229_n400# a_29_n497# a_n29_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LUSSBJ a_108_n288# a_50_n200# a_n208_n288# a_n400_n422#
+ a_n108_n200# a_n266_n200# a_n50_n288# a_208_n200#
X0 a_n108_n200# a_n208_n288# a_n266_n200# a_n400_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_208_n200# a_108_n288# a_50_n200# a_n400_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_50_n200# a_n50_n288# a_n108_n200# a_n400_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__res_high_po_2p85_EP2UD7 a_n2283_n3624# a_381_n3624# a_n2437_n3778#
+ a_n285_3192# a_1047_3192# a_n951_3192# a_1713_3192# a_n1617_n3624# a_381_3192# a_n285_n3624#
+ a_n951_n3624# a_1047_n3624# a_n2283_3192# a_1713_n3624# a_n1617_3192#
X0 a_n285_3192# a_n285_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X1 a_1047_3192# a_1047_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X2 a_n951_3192# a_n951_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X3 a_1713_3192# a_1713_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X4 a_n2283_3192# a_n2283_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X5 a_n1617_3192# a_n1617_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X6 a_381_3192# a_381_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HHHAEV a_n29_n400# a_n229_n488# a_n421_n622#
+ a_n287_n400# a_229_n400# a_29_n488#
X0 a_229_n400# a_29_n488# a_n29_n400# a_n421_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X1 a_n29_n400# a_n229_n488# a_n287_n400# a_n421_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TAUUP3 a_n345_n431# a_129_n431# a_29_n457# a_n129_n457#
+ a_287_n431# a_187_n457# a_n287_n457# a_n29_n431# a_n479_n591# a_n187_n431#
X0 a_n187_n431# a_n287_n457# a_n345_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_287_n431# a_187_n457# a_129_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_129_n431# a_29_n457# a_n29_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n29_n431# a_n129_n457# a_n187_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RJSTGP a_29_n297# a_n887_n200# a_n29_n200# a_n829_n297#
+ w_n1087_n497# a_829_n200#
X0 a_n29_n200# a_n829_n297# a_n887_n200# w_n1087_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=4
X1 a_829_n200# a_29_n297# a_n29_n200# w_n1087_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8JQF8T a_n100_n1015# a_n158_118# a_n100_21# w_n358_n1215#
+ a_100_n918# a_n158_n918# a_100_118#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n1215# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X1 a_100_n918# a_n100_n1015# a_n158_n918# w_n358_n1215# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PNRDLC a_n150_n897# a_150_n800# w_n408_n1097#
+ a_n208_n800#
X0 a_150_n800# a_n150_n897# a_n208_n800# w_n408_n1097# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_46Z5PG a_129_n200# a_29_n288# a_n129_n288# a_n321_n422#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RRA4TL a_n258_n50# a_n200_n138# a_200_n50# a_n392_n272#
X0 a_200_n50# a_n200_n138# a_n258_n50# a_n392_n272# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CRL9SD a_n150_n897# a_150_n800# w_n408_n1097#
+ a_n208_n800#
X0 a_150_n800# a_n150_n897# a_n208_n800# w_n408_n1097# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__pfet_01v8_YTEHH6 w_n425_n619# a_n29_n400# a_29_n497# a_n287_n400#
+ a_n229_n497# a_229_n400#
X0 a_n29_n400# a_n229_n497# a_n287_n400# w_n425_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_229_n400# a_29_n497# a_n29_n400# w_n425_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_8TUSME a_n345_n200# a_129_n200# a_287_n200# a_n479_n422#
+ a_29_n288# a_n129_n288# a_187_n288# a_n287_n288# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n288# a_n29_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n288# a_n187_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T8W2FW a_150_n800# a_n208_n800# a_n150_n888#
+ a_n342_n1022#
X0 a_150_n800# a_n150_n888# a_n208_n800# a_n342_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_AUB4P8 a_150_n800# a_n208_n800# a_n150_n888#
+ a_n342_n1022#
X0 a_150_n800# a_n150_n888# a_n208_n800# a_n342_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__nfet_01v8_HWT53N a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_EPRAC4 a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LHNF5N a_n345_n431# a_129_n431# a_29_n457# a_n129_n457#
+ a_287_n431# a_187_n457# a_n287_n457# a_n29_n431# a_n479_n591# a_n187_n431#
X0 a_n187_n431# a_n287_n457# a_n345_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_287_n431# a_187_n457# a_129_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_129_n431# a_29_n457# a_n29_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n29_n431# a_n129_n457# a_n187_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Q8UPKT a_n829_n615# w_n1087_n815# a_29_n615#
+ a_29_21# a_n887_n518# a_829_118# a_n29_n518# a_829_n518# a_n29_118# a_n887_118#
+ a_n829_21#
X0 a_829_n518# a_29_n615# a_n29_n518# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=4
X1 a_829_118# a_29_21# a_n29_118# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=4
X2 a_n29_118# a_n829_21# a_n887_118# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=4
X3 a_n29_n518# a_n829_n615# a_n887_n518# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_X332GA a_29_n297# a_n129_n297# a_129_n200# a_n29_n200#
+ w_n387_n497# a_n187_n200#
X0 a_129_n200# a_29_n297# a_n29_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n297# a_n187_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_4RA4DJ a_n603_n288# a_n345_n200# a_129_n200#
+ a_n503_n200# a_287_n200# a_n661_n200# a_445_n200# a_29_n288# a_n129_n288# a_603_n200#
+ a_187_n288# a_n795_n422# a_n287_n288# a_345_n288# a_n29_n200# a_n187_n200# a_n445_n288#
+ a_503_n288#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n288# a_n503_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_129_n200# a_29_n288# a_n29_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n288# a_287_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n503_n200# a_n603_n288# a_n661_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X6 a_n29_n200# a_n129_n288# a_n187_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X7 a_603_n200# a_503_n288# a_445_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_GHE6BF a_n158_n518# a_n158_118# a_n100_21# a_n100_n615#
+ w_n358_n815# a_100_118# a_100_n518#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_n518# a_n100_n615# a_n158_n518# w_n358_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WGHV7X a_400_n509# a_n458_109# a_n400_21# a_n458_n509#
+ a_n592_n731# a_400_109# a_n400_n597#
X0 a_400_n509# a_n400_n597# a_n458_n509# a_n592_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X1 a_400_109# a_n400_21# a_n458_109# a_n592_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LURNA9 a_n287_n200# a_n1061_n200# a_745_n200#
+ a_n487_n288# a_545_n288# a_229_n200# a_n1195_n422# a_n545_n200# a_29_n288# a_n745_n288#
+ a_1003_n200# a_803_n288# a_487_n200# a_n29_n200# a_n229_n288# a_287_n288# a_n1003_n288#
+ a_n803_n200#
X0 a_487_n200# a_287_n288# a_229_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n288# a_n287_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_229_n200# a_29_n288# a_n29_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n545_n200# a_n745_n288# a_n803_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n803_n200# a_n1003_n288# a_n1061_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X5 a_n287_n200# a_n487_n288# a_n545_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_745_n200# a_545_n288# a_487_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_1003_n200# a_803_n288# a_745_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RM8L2M a_n258_n50# a_n200_n138# a_200_n50# a_n392_n272#
X0 a_200_n50# a_n200_n138# a_n258_n50# a_n392_n272# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HDHSEV a_n29_n400# a_n229_n488# a_n421_n622#
+ a_n287_n400# a_229_n400# a_29_n488#
X0 a_229_n400# a_29_n488# a_n29_n400# a_n421_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X1 a_n29_n400# a_n229_n488# a_n287_n400# a_n421_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_N8ANR9 a_n345_n364# a_129_n364# a_287_n364# w_n545_n662#
+ a_29_n461# a_n129_n461# a_187_n461# a_n287_n461# a_n29_n364# a_n187_n364#
X0 a_n187_n364# a_n287_n461# a_n345_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_287_n364# a_187_n461# a_129_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_129_n364# a_29_n461# a_n29_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n29_n364# a_n129_n461# a_n187_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6UJQA2 a_n187_n436# a_n345_n436# a_129_n436#
+ a_287_n436# w_n545_n662# a_29_n462# a_n129_n462# a_187_n462# a_n287_n462# a_n29_n436#
X0 a_129_n436# a_29_n462# a_n29_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n436# a_n129_n462# a_n187_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_n187_n436# a_n287_n462# a_n345_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X3 a_287_n436# a_187_n462# a_129_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CDNABP a_n100_n597# a_n100_21# a_100_109# a_100_n509#
+ a_n158_n509# a_n292_n731# a_n158_109#
X0 a_100_n509# a_n100_n597# a_n158_n509# a_n292_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_109# a_n100_21# a_n158_109# a_n292_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CS979Q a_n400_n615# a_400_118# w_n658_n815# a_n400_21#
+ a_400_n518# a_n458_118# a_n458_n518#
X0 a_400_118# a_n400_21# a_n458_118# w_n658_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X1 a_400_n518# a_n400_n615# a_n458_n518# w_n658_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_2CKAKF a_n819_n200# a_n345_n200# a_n977_n200#
+ a_n1135_n200# a_29_n297# a_n129_n297# a_187_n297# a_129_n200# a_n503_n200# a_n1293_n200#
+ a_n287_n297# a_819_n297# a_345_n297# a_n1077_n297# a_287_n200# a_n661_n200# a_n919_n297#
+ a_977_n297# a_n445_n297# a_919_n200# a_503_n297# a_n1235_n297# a_445_n200# a_1135_n297#
+ a_n603_n297# a_1077_n200# a_661_n297# a_603_n200# w_n1493_n497# a_n761_n297# a_1235_n200#
+ a_761_n200# a_n29_n200# a_n187_n200#
X0 a_n819_n200# a_n919_n297# a_n977_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n661_n200# a_n761_n297# a_n819_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_919_n200# a_819_n297# a_761_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n187_n200# a_n287_n297# a_n345_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_761_n200# a_661_n297# a_603_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X5 a_287_n200# a_187_n297# a_129_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X6 a_n345_n200# a_n445_n297# a_n503_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X7 a_129_n200# a_29_n297# a_n29_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X8 a_445_n200# a_345_n297# a_287_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X9 a_n977_n200# a_n1077_n297# a_n1135_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X10 a_n503_n200# a_n603_n297# a_n661_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X11 a_1077_n200# a_977_n297# a_919_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X12 a_n29_n200# a_n129_n297# a_n187_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X13 a_603_n200# a_503_n297# a_445_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X14 a_n1135_n200# a_n1235_n297# a_n1293_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X15 a_1235_n200# a_1135_n297# a_1077_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EEFBWQ a_400_n200# a_n592_n422# a_n458_n200#
+ a_n400_n288#
X0 a_400_n200# a_n400_n288# a_n458_n200# a_n592_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_9432CF a_n345_n200# a_29_n297# a_n129_n297# w_n703_n497#
+ a_187_n297# a_129_n200# a_n503_n200# a_n287_n297# a_345_n297# a_287_n200# a_n445_n297#
+ a_445_n200# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n297# a_129_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n297# a_n503_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_129_n200# a_29_n297# a_n29_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n297# a_287_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n29_n200# a_n129_n297# a_n187_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_2432J2 a_n345_n200# a_29_n297# a_n129_n297# a_187_n297#
+ a_129_n200# a_n287_n297# a_287_n200# a_n29_n200# a_n187_n200# w_n545_n497#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n297# a_129_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n297# a_n29_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n297# a_n187_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_ak_ip__comparator Vinp Vinm AVDD AGND en hyst[1] hyst[0] trim[5] trim[4]
+ trim[3] trim[2] trim[1] trim[0] Vout DVDD ibias DGND
Xlevel_shifter_up_3 AVDD en en_hv enb_hv DVDD DGND m1_36128_n32592# AGND level_shifter_up
Xsky130_fd_pr__pfet_g5v0d10v5_RUG6CB_0 m1_25710_11400# AVDD AVDD m1_25710_11400# sky130_fd_pr__pfet_g5v0d10v5_RUG6CB
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_82 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_60 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_REE66T_1 m1_36250_n26840# m1_2500_n30560# m1_2500_n30560#
+ m1_36250_n26840# m1_31820_n13600# m1_36250_n26840# m1_31820_n13600# m1_2500_n30560#
+ m1_36250_n26840# m1_36250_n26840# m1_31820_n13600# m1_36250_n26840# m1_36250_n26840#
+ m1_36250_n26840# m1_31820_n13600# m1_2500_n30560# AVDD m1_2500_n30560# sky130_fd_pr__pfet_g5v0d10v5_REE66T
Xlevel_shifter_up_4 AVDD trim[3] level_shifter_up_4/x_hv trim3b_hv DVDD DGND m1_35128_n32592#
+ AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_LUSSBJ_0 hyst0_hv AGND hyst0_hv AGND m1_33660_n1540#
+ AGND hyst0_hv m1_33660_n1540# sky130_fd_pr__nfet_g5v0d10v5_LUSSBJ
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_61 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_83 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_50 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__res_high_po_2p85_EP2UD7_0 AGND m1_25040_4590# AGND m1_24380_11400#
+ m1_25710_11400# m1_23050_11400# AGND m1_23040_4590# m1_24380_11400# m1_23710_4590#
+ m1_23710_4590# m1_25040_4590# AGND AGND m1_23050_11400# sky130_fd_pr__res_high_po_2p85_EP2UD7
Xlevel_shifter_up_5 AVDD trim[4] level_shifter_up_5/x_hv trim4b_hv DVDD DGND m1_34128_n32592#
+ AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_40 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_73 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_84 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_62 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_51 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__res_high_po_2p85_EP2UD7_1 AGND m1_24360_n31900# AGND m1_23690_n25080#
+ m1_25020_n25080# m1_23690_n25080# AGND m1_23030_n31900# m1_25020_n25080# m1_24360_n31900#
+ m1_23030_n31900# res_p_bot AGND AGND m1_23030_n25080# sky130_fd_pr__res_high_po_2p85_EP2UD7
Xlevel_shifter_up_6 AVDD trim[0] level_shifter_up_6/x_hv level_shifter_up_6/xb_hv
+ DVDD DGND level_shifter_up_6/m1_380_440# AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_74 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_85 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_63 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_41 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_30 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_52 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xlevel_shifter_up_7 AVDD trim[2] level_shifter_up_7/x_hv level_shifter_up_7/xb_hv
+ DVDD DGND level_shifter_up_7/m1_380_440# AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_53 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_31 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_75 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_42 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_20 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_86 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xlevel_shifter_up_8 AVDD trim[1] level_shifter_up_8/x_hv level_shifter_up_8/xb_hv
+ DVDD DGND level_shifter_up_8/m1_380_440# AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_32 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_76 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_54 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_43 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_21 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_87 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_10 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_HHHAEV_0 DGND m1_30900_4740# DGND m1_35900_10510# m1_30900_4740#
+ m1_30900_4740# sky130_fd_pr__nfet_g5v0d10v5_HHHAEV
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_77 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_55 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_33 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_22 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_88 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_11 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_44 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_78 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_23 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_34 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_12 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_TAUUP3_0 bias_n AGND enb_hv enb_hv bias_n enb_hv enb_hv
+ bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5_TAUUP3
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_45 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_RJSTGP_0 m1_29940_7140# AVDD m1_29940_7140# m1_29940_7140#
+ AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_RJSTGP
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_79 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_57 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_35 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_13 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_8JQF8T_0 Vop m1_29860_5120# Vom AVDD m1_29880_4800#
+ m1_29860_5120# m1_30900_4740# sky130_fd_pr__pfet_g5v0d10v5_8JQF8T
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_46 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_14 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_58 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_36 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_30 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_25 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_46Z5PG_0 AGND level_shifter_up_8/x_hv level_shifter_up_8/x_hv
+ AGND m1_32060_2060# AGND sky130_fd_pr__nfet_g5v0d10v5_46Z5PG
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_15 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_59 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_37 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_31 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_20 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_26 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_RRA4TL_0 m1_29880_4800# m1_30900_4740# DGND DGND sky130_fd_pr__nfet_g5v0d10v5_RRA4TL
Xsky130_fd_pr__nfet_g5v0d10v5_46Z5PG_1 AGND level_shifter_up_6/x_hv level_shifter_up_6/x_hv
+ AGND m1_35270_2060# AGND sky130_fd_pr__nfet_g5v0d10v5_46Z5PG
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_49 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_38 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_32 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|2] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|2] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|2] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|2] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|3] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|3] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|3] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|3] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|4] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|4] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|4] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|4] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|5] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|5] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|5] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|5] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_21 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_10 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_27 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_01v8_YTEHH6_0 DVDD m1_35390_11200# m1_35390_11200# DVDD m1_35390_11200#
+ DVDD sky130_fd_pr__pfet_01v8_YTEHH6
Xsky130_fd_pr__nfet_g5v0d10v5_8TUSME_0 DGND m1_35900_10510# DGND DGND enb_hv enb_hv
+ enb_hv enb_hv DGND m1_35900_10510# sky130_fd_pr__nfet_g5v0d10v5_8TUSME
Xsky130_fd_pr__nfet_g5v0d10v5_46Z5PG_2 AGND level_shifter_up_8/x_hv level_shifter_up_8/x_hv
+ AGND m1_32060_2060# AGND sky130_fd_pr__nfet_g5v0d10v5_46Z5PG
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_28 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_33 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_22 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_11 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_17 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_01v8_YTEHH6_1 DVDD m1_35900_10510# m1_35390_11200# DVDD m1_35390_11200#
+ DVDD sky130_fd_pr__pfet_01v8_YTEHH6
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_30 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_29 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_34 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_23 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_12 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_AUB4P8_0 m1_9080_4100# m1_7790_4530# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_AUB4P8
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_18 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_31 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_20 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_01v8_HWT53N_0 DGND m1_35900_10510# m1_34800_n26840# DGND sky130_fd_pr__nfet_01v8_HWT53N
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_35 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_24 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_13 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_AUB4P8_1 m1_9080_4100# m1_7790_4530# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_AUB4P8
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_19 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_32 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_21 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_10 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_01v8_HWT53N_1 DGND m1_36250_n26840# Vout DGND sky130_fd_pr__nfet_01v8_HWT53N
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_9 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_01v8_EPRAC4_0 Vout DVDD m1_36250_n26840# DVDD sky130_fd_pr__pfet_01v8_EPRAC4
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_25 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_14 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_0 m1_23030_n25080# m1_4100_n29230# trim5b_hv
+ trim5b_hv m1_23030_n25080# trim5b_hv trim5b_hv m1_23030_n25080# AGND m1_4100_n29230#
+ sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_33 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_22 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_11 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_01v8_HWT53N_2 DGND m1_34800_n26840# m1_36250_n26840# DGND sky130_fd_pr__nfet_01v8_HWT53N
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_26 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_15 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_01v8_EPRAC4_1 m1_34800_n26840# DVDD m1_35900_10510# DVDD sky130_fd_pr__pfet_01v8_EPRAC4
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_1 res_p_bot m1_4100_n28430# trim5b_hv trim5b_hv
+ res_p_bot trim5b_hv trim5b_hv res_p_bot AGND m1_4100_n28430# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_34 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_23 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_12 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_01v8_EPRAC4_2 m1_36250_n26840# DVDD m1_34800_n26840# DVDD sky130_fd_pr__pfet_01v8_EPRAC4
Xsky130_fd_pr__pfet_g5v0d10v5_Q8UPKT_0 m1_29940_7140# AVDD m1_29940_7140# m1_29940_7140#
+ AVDD AVDD m1_29860_5120# AVDD m1_29860_5120# AVDD m1_29940_7140# sky130_fd_pr__pfet_g5v0d10v5_Q8UPKT
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_27 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_16 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_2 m1_23030_n25080# m1_4100_n28430# trim5_hv trim5_hv
+ m1_23030_n25080# trim5_hv trim5_hv m1_23030_n25080# AGND m1_4100_n28430# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_35 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_24 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_17 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_28 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_3 m1_27260_n27254# m1_23030_n25080# trim3b_hv
+ trim3b_hv m1_27260_n27254# trim3b_hv trim3b_hv m1_27260_n27254# AGND m1_23030_n25080#
+ sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_25 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_29 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_18 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_4 res_p_bot m1_4100_n29230# trim5_hv trim5_hv
+ res_p_bot trim5_hv trim5_hv res_p_bot AGND m1_4100_n29230# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_26 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_15 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_19 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_5 res_p_bot m1_27260_n27254# trim4b_hv trim4b_hv
+ res_p_bot trim4b_hv trim4b_hv res_p_bot AGND m1_27260_n27254# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_27 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_16 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_X332GA_0 trim3b_hv trim3b_hv AVDD m1_33660_n22250# AVDD
+ AVDD sky130_fd_pr__pfet_g5v0d10v5_X332GA
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_17 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_4RA4DJ_0 hyst1_hv AGND m1_32060_n3340# m1_32060_n3340#
+ AGND AGND m1_32060_n3340# hyst1_hv hyst1_hv AGND hyst1_hv AGND hyst1_hv hyst1_hv
+ AGND m1_32060_n3340# hyst1_hv hyst1_hv sky130_fd_pr__nfet_g5v0d10v5_4RA4DJ
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_28 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|0] res_p_bot res_p_bot casc_p casc_p AVDD
+ m1_11260_n21330# m1_11260_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|0] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|0] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|0] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|0] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|0] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|1] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|1] m1_12400_n19010# m1_12400_n19010# casc_p
+ casc_p AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|1] m1_12400_n19010# m1_12400_n19010# casc_p
+ casc_p AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|1] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|1] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|1] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|2] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|2] bias_var_n bias_var_n casc_p casc_p AVDD
+ m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|2] bias_var_n bias_var_n casc_p casc_p AVDD
+ m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|2] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|2] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|2] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|3] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|3] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|3] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|3] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|3] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|3] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|4] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|4] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|4] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|4] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|4] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|4] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|5] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|5] m1_12860_n11800# m1_12860_n11800# casc_p
+ casc_p AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|5] m1_12860_n11800# m1_12860_n11800# casc_p
+ casc_p AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|5] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|5] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|5] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|6] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|6] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|6] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|6] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|6] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|6] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|7] m1_11180_n8390# m1_11180_n8390# m1_11180_n8390#
+ m1_11180_n8390# AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|7] m1_11180_n8390# m1_11180_n8390# m1_11180_n8390#
+ m1_11180_n8390# AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|7] m1_11180_n8390# m1_11180_n8390# m1_11180_n8390#
+ m1_11180_n8390# AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|7] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|7] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|7] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|0] m1_11260_n4491# AGND bias_n AGND AGND
+ m1_11260_n4491# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|0] m1_12840_n4260# AGND bias_n m1_12600_n4860#
+ AGND m1_12840_n4260# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|0] m1_14440_n4260# AGND bias_n m1_14200_n4860#
+ AGND m1_14440_n4260# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|0] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|0] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|0] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|0] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|0] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|0] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|0] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|0] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|0] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|1] m1_11260_n2671# AGND bias_n AGND AGND
+ m1_11260_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|1] m1_12860_n2671# AGND bias_n AGND AGND
+ m1_12860_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|1] m1_14459_n2671# AGND bias_n AGND AGND
+ m1_14459_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|1] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|1] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|1] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|1] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|1] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|1] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|1] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|1] m1_33659_n2671# m1_33660_n1540# bias_n
+ m1_33660_n1540# AGND m1_33659_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|1] m1_33659_n2671# AGND AGND m1_33660_n1540#
+ AGND AGND bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|2] bias_n AGND bias_n AGND AGND bias_n bias_n
+ sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|2] casc_n AGND bias_n AGND AGND casc_n bias_n
+ sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|2] bias_var_n AGND bias_var_n AGND AGND bias_var_n
+ bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|2] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|2] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|2] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|2] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|2] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|2] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|2] m1_32060_n890# AGND m1_12400_n19010#
+ AGND AGND m1_32060_n890# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|2] m1_32060_n890# AGND m1_12400_n19010#
+ AGND AGND m1_32060_n890# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|2] m1_32060_n890# AGND m1_12400_n19010#
+ AGND AGND m1_32060_n890# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|3] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|3] bias_n m1_11240_2060# ibias m1_11240_2060#
+ AGND m1_11860_1120# ibias sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|3] m1_11860_1120# m1_12840_2060# ibias m1_12840_2060#
+ AGND ibias ibias sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|3] m1_12400_n19010# AGND m1_12400_n19010#
+ AGND AGND m1_12400_n19010# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|3] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|3] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|3] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|3] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|3] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|3] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|3] m1_32060_910# m1_32060_2060# bias_n m1_32060_2060#
+ AGND m1_32060_910# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|3] m1_32060_910# m1_32060_2060# bias_n m1_32060_2060#
+ AGND m1_32060_910# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|3] m1_35259_929# m1_35270_2060# bias_n m1_35270_2060#
+ AGND m1_35259_929# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|3] m1_36870_930# AGND bias_n AGND AGND m1_37480_930#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_29 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_18 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_0 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_19 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_1 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_2 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_0 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_3 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_1 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_4 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_2 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LURNA9_0 m1_32060_n4840# m1_2500_5340# m1_32060_n4840#
+ m1_34800_n26840# m1_34800_n26840# m1_32060_n4840# AGND m1_2500_5340# m1_34800_n26840#
+ m1_34800_n26840# m1_2500_5340# m1_34800_n26840# m1_2500_5340# m1_2500_5340# m1_34800_n26840#
+ m1_34800_n26840# m1_34800_n26840# m1_32060_n4840# sky130_fd_pr__nfet_g5v0d10v5_LURNA9
Xsky130_fd_pr__nfet_g5v0d10v5_RM8L2M_0 DGND m1_29880_4800# m1_30900_4740# DGND sky130_fd_pr__nfet_g5v0d10v5_RM8L2M
Xsky130_fd_pr__nfet_g5v0d10v5_HDHSEV_0 DGND m1_29880_4800# DGND m1_35390_11200# m1_29880_4800#
+ m1_29880_4800# sky130_fd_pr__nfet_g5v0d10v5_HDHSEV
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_5 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_0 m1_23040_4590# m1_4100_9160# m1_23040_4590#
+ AVDD level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv
+ level_shifter_up_7/xb_hv m1_23040_4590# m1_4100_9160# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_3 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LURNA9_1 m1_32060_n4840# m1_2500_6140# m1_32060_n4840#
+ m1_36250_n26840# m1_36250_n26840# m1_32060_n4840# AGND m1_2500_6140# m1_36250_n26840#
+ m1_36250_n26840# m1_2500_6140# m1_36250_n26840# m1_2500_6140# m1_2500_6140# m1_36250_n26840#
+ m1_36250_n26840# m1_36250_n26840# m1_32060_n4840# sky130_fd_pr__nfet_g5v0d10v5_LURNA9
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_1 m1_25710_11400# m1_27260_9746# m1_25710_11400#
+ AVDD level_shifter_up_6/x_hv level_shifter_up_6/x_hv level_shifter_up_6/x_hv level_shifter_up_6/x_hv
+ m1_25710_11400# m1_27260_9746# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_6UJQA2_0 AVDD bias_p AVDD bias_p AVDD en_hv en_hv en_hv
+ en_hv bias_p sky130_fd_pr__pfet_g5v0d10v5_6UJQA2
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|0] casc_n casc_n casc_p casc_p m1_11260_n4491#
+ AGND m1_11260_n4491# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|0] casc_n casc_n m1_11180_n8390# m1_12600_n4860#
+ m1_12850_n4460# AGND m1_12850_n4460# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|0] casc_n casc_n m1_12860_n11800# m1_14200_n4860#
+ m1_14450_n4460# AGND m1_14450_n4460# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|0] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|0] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|0] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|1] casc_n casc_n bias_p bias_p m1_11260_n2671#
+ AGND m1_11260_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|1] casc_n casc_n m1_9080_4100# m1_9080_4100#
+ m1_12860_n2671# AGND m1_12860_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|1] casc_n casc_n m1_2120_n22080# m1_2120_n22080#
+ m1_14459_n2671# AGND m1_14459_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|1] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|1] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_33659_n2671# AGND m1_33659_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|1] casc_n casc_n casc_n m1_32060_n4840#
+ m1_33659_n2671# AGND casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|2] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|2] ibias ibias AVDD AVDD casc_n AGND casc_n
+ sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|2] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|2] casc_n casc_n m1_420_6500# m1_420_6500#
+ m1_32060_n890# AGND m1_32060_n890# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|2] casc_n casc_n m1_420_6500# m1_420_6500#
+ m1_32060_n890# AGND m1_32060_n890# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|2] casc_n casc_n m1_420_6500# m1_420_6500#
+ m1_32060_n890# AGND m1_32060_n890# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|3] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|3] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|3] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|3] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|3] casc_n casc_n m1_23040_4590# m1_23040_4590#
+ m1_32060_910# AGND m1_32060_910# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|3] casc_n casc_n m1_23040_4590# m1_23040_4590#
+ m1_32060_910# AGND m1_32060_910# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|3] casc_n casc_n m1_23040_4590# m1_23040_4590#
+ m1_35259_929# AGND m1_35259_929# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|3] casc_n casc_n m1_29940_7140# m1_25710_11400#
+ m1_36870_930# AGND m1_37480_930# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_6 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_4 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_2 m1_27260_9746# m1_23040_4590# m1_27260_9746#
+ AVDD level_shifter_up_8/x_hv level_shifter_up_8/x_hv level_shifter_up_8/x_hv level_shifter_up_8/x_hv
+ m1_27260_9746# m1_23040_4590# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_5 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|0] bias_p AVDD AVDD bias_p AVDD m1_11260_n21330#
+ m1_11260_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|0] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|0] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|0] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|0] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|0] bias_p m1_33660_n22250# AVDD bias_p m1_33660_n22250#
+ m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|0] bias_p m1_33660_n22250# AVDD bias_p m1_33660_n22250#
+ m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|1] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|1] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|1] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|1] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|1] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|1] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|2] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|2] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|2] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|3] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|3] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|3] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|4] bias_p AVDD AVDD bias_p AVDD m1_11260_n14130#
+ m1_11260_n14130# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|4] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|4] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|4] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|4] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|4] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|4] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|5] bias_p m1_11260_n14130# AVDD bias_p m1_11260_n14130#
+ m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|5] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|5] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|5] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|5] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|5] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|5] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|6] bias_p AVDD AVDD bias_p AVDD bias_p bias_p
+ sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|6] bias_p AVDD AVDD bias_p AVDD bias_p bias_p
+ sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|6] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|6] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|6] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|6] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|6] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|6] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|7] m1_11180_n8390# AVDD AVDD m1_11180_n8390#
+ AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|7] casc_p m1_11260_n8730# AVDD casc_p m1_11260_n8730#
+ casc_p casc_p sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|7] casc_p m1_11260_n8730# AVDD casc_p m1_11260_n8730#
+ casc_p casc_p sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|7] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|7] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|7] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|7] bias_p m1_32060_n9640# AVDD bias_p m1_32060_n9640#
+ m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|7] bias_p m1_32060_n9640# AVDD bias_p m1_32060_n9640#
+ m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|7] bias_p m1_32060_n9640# AVDD bias_p m1_32060_n9640#
+ m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_7 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_2CKAKF_0 m1_32060_n15040# AVDD AVDD m1_32060_n15040#
+ hyst1b_hv hyst1b_hv hyst1b_hv m1_32060_n15040# m1_32060_n15040# AVDD hyst1b_hv hyst1b_hv
+ hyst1b_hv hyst1b_hv AVDD AVDD hyst1b_hv hyst1b_hv hyst1b_hv AVDD hyst1b_hv hyst1b_hv
+ m1_32060_n15040# hyst1b_hv hyst1b_hv m1_32060_n15040# hyst1b_hv AVDD AVDD hyst1b_hv
+ AVDD m1_32060_n15040# AVDD m1_32060_n15040# sky130_fd_pr__pfet_g5v0d10v5_2CKAKF
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_8 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_3 m1_25710_11400# m1_4100_9160# m1_25710_11400#
+ AVDD level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv
+ m1_25710_11400# m1_4100_9160# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_6 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_EEFBWQ_0 AGND AGND res_p_bot res_p_bot sky130_fd_pr__nfet_g5v0d10v5_EEFBWQ
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_4 m1_25710_11400# m1_4100_8360# m1_25710_11400#
+ AVDD level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv
+ level_shifter_up_7/xb_hv m1_25710_11400# m1_4100_8360# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_7 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_9 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xlevel_shifter_up_0 AVDD trim[5] trim5_hv trim5b_hv DVDD DGND m1_33128_n32592# AGND
+ level_shifter_up
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_5 m1_23040_4590# m1_4100_8360# m1_23040_4590#
+ AVDD level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv
+ m1_23040_4590# m1_4100_8360# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_8 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_9432CF_0 AVDD hyst0b_hv hyst0b_hv AVDD hyst0b_hv m1_32060_n9640#
+ m1_32060_n9640# hyst0b_hv hyst0b_hv AVDD hyst0b_hv m1_32060_n9640# AVDD m1_32060_n9640#
+ sky130_fd_pr__pfet_g5v0d10v5_9432CF
Xlevel_shifter_up_1 AVDD level_shifter_up_1/x_lv hyst0_hv hyst0b_hv DVDD DGND m1_38128_n32592#
+ AGND level_shifter_up
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_9 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xlevel_shifter_up_2 AVDD level_shifter_up_2/x_lv hyst1_hv hyst1b_hv DVDD DGND m1_37128_n32592#
+ AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_81 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_2432J2_1 AVDD trim4b_hv trim4b_hv trim4b_hv m1_32060_n22250#
+ trim4b_hv AVDD AVDD m1_32060_n22250# AVDD sky130_fd_pr__pfet_g5v0d10v5_2432J2
Xsky130_fd_pr__pfet_g5v0d10v5_REE66T_0 m1_34800_n26840# Vfold_bot_m Vfold_bot_m m1_34800_n26840#
+ m1_31820_n13600# m1_34800_n26840# m1_31820_n13600# Vfold_bot_m m1_34800_n26840#
+ m1_34800_n26840# m1_31820_n13600# m1_34800_n26840# m1_34800_n26840# m1_34800_n26840#
+ m1_31820_n13600# Vfold_bot_m AVDD Vfold_bot_m sky130_fd_pr__pfet_g5v0d10v5_REE66T
.ends

.subckt lpopamp_slice im ip o en enb avdd avss bpa bpb bnb bna xp ypm ypp zpm zpp
+ xn ynm ynp znm znp vsub
X0 a_38000_1800# znp a_37700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1 o znm a_71000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X3 a_75200_n3300# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X4 a_34700_1800# znp a_34400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X5 ynp znp a_53600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X6 o znm a_73400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X7 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X8 ypp zpp a_45800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X9 a_31400_1800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X10 a_57800_n3300# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X11 a_70400_1800# znp a_70100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X12 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X13 a_20300_n3300# bna a_20000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X14 a_24200_n3300# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X15 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X16 a_73400_n1600# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X17 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X18 znp znp a_51800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X19 a_56000_n1600# znp a_55700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X20 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X21 a_31400_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X22 a_63200_10000# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X23 ynm znp a_59600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X24 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X25 a_70400_6100# zpp a_70100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X26 a_27200_7400# zpp a_26900_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X27 ypp zpp a_41600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X28 a_22400_n1600# bna a_22100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X29 ynm znp a_59600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X30 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X31 a_45800_10000# zpp a_45500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X32 xn im a_26000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X33 a_17600_1800# bna a_17300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X34 a_49700_10000# bpa a_49400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X35 a_56600_1800# znp a_56300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X36 a_29000_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X37 bna_ bnb a_14000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X38 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X39 a_51800_100# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X40 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X41 znp znp a_53000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X42 a_25700_8700# zpp a_25400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X43 a_64700_8700# zpp a_64400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X44 a_22400_8700# zpp a_22100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X45 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X46 a_8600_1800# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X47 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X48 znm bnb a_63800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X49 a_68000_n3300# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X50 a_44000_100# bnb a_43700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X51 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X52 bnb bnb a_5000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X53 a_17600_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X54 a_200_n3300# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X55 a_30500_n3300# bna a_30200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X56 a_11000_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X57 a_56600_6100# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X58 a_34400_n3300# znp a_34100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X59 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X60 znp znp a_53000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X61 avdd bpa a_53000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X62 bna_ bnb a_12800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X63 ynm znp a_38000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X64 a_17000_n3300# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X65 a_20300_100# bna a_20000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X66 a_16100_7400# bpa a_15800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X67 a_39500_1800# znp a_39200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X68 a_55100_7400# bpb a_54800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X69 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X70 a_8600_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X71 a_36200_1800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X72 a_51800_7400# bpb a_51500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X73 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X74 a_70100_n1600# znp a_69800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X75 bnb bnb a_3800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X76 a_45500_100# bnb a_45200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X77 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X78 a_75200_1800# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X79 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X80 a_8000_n3300# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X81 wp bpb a_51800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X82 a_32600_n1600# znp a_32300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X83 a_1400_100# bna a_1100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X84 bnb bnb a_12200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X85 a_56000_10000# bpb a_55700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X86 a_36500_n1600# znp a_36200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X87 a_44300_8700# zpp a_44000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X88 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X89 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X90 a_22400_10000# zpp a_22100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X91 bpb bna a_18800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X92 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X93 avdd zpp a_26000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X94 a_37700_100# znp a_37400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X95 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X96 a_36200_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X97 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X98 bnb bnb a_9800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X99 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X100 avss znp a_40400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X101 a_29900_100# bna a_29600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X102 a_44600_n3300# bnb a_44300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X103 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X104 a_48500_n3300# bna a_48200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X105 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X106 a_31400_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X107 a_39200_100# znp a_38900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X108 xn im a_24800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X109 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X110 a_27200_8700# zpp a_26900_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X111 znm bnb a_63800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X112 a_70400_7400# zpp a_70100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X113 a_21800_1800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X114 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X115 a_60800_1800# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X116 a_60200_n1600# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X117 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X118 a_42800_n1600# bna a_42500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X119 wn bnb a_46400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X120 a_70100_10000# zpp a_69800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X121 ypp zpp a_24800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X122 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X123 avdd zpp a_63800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X124 a_36500_10000# bpa a_36200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X125 a_21800_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X126 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X127 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X128 a_17600_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X129 avdd bpa a_18800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X130 a_56600_7400# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X131 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X132 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X133 a_47000_1800# bna wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X134 avdd bpa a_53000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X135 znm znp a_60200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X136 a_72200_n3300# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X137 a_50900_n3300# znp a_50600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X138 a_43700_1800# bnb a_43400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X139 a_16100_8700# bpa a_15800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X140 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X141 a_54800_n3300# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X142 a_55100_8700# bpb a_54800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X143 a_40400_1800# znp a_40100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X144 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X145 a_58700_n3300# znp a_58400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X146 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X147 a_8600_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X148 a_51800_8700# bpb a_51500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X149 a_21200_n3300# bna a_20900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X150 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X151 ynp znp a_52400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X152 a_70400_n1600# znp a_70100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X153 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X154 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X155 avss znm a_74000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X156 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X157 a_53000_n1600# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X158 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X159 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X160 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X161 a_56900_n1600# znp a_56600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X162 a_40400_6100# bpa a_40100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X163 zpp bnb a_44600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X164 a_36200_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X165 a_29900_1800# bna a_29600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X166 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X167 a_23300_n1600# bna a_23000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X168 bna_ bnb a_11600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X169 a_68900_1800# znp a_68600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X170 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X171 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X172 a_27200_n1600# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X173 a_26600_1800# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X174 a_54200_100# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X175 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X176 a_70100_100# znp a_69800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X177 a_65600_1800# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X178 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X179 a_23300_1800# bna a_23000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X180 a_21200_100# bna a_20900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X181 a_37100_100# znp a_36800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X182 zpm bnb a_62000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X183 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X184 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X185 a_31400_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X186 a_70400_8700# zpp a_70100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X187 ynm znp a_60800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X188 a_46400_100# bnb a_46100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X189 ypm zpp a_29600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X190 a_65000_n3300# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X191 bna_ bna a_2000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X192 a_13400_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X193 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X194 a_68900_n3300# znp a_68600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X195 a_26600_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X196 a_31400_n3300# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X197 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X198 a_23300_6100# zpp a_23000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X199 a_35300_n3300# znp a_35000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X200 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X201 a_14000_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X202 a_39200_n3300# znp a_38900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X203 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X204 a_38600_100# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X205 a_17900_n3300# bna a_17600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X206 ypp zpp a_24800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X207 a_48500_1800# bna a_48200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X208 avdd zpp a_63800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X209 a_21800_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X210 a_70400_10000# zpp a_70100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X211 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X212 ynm znp a_66800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X213 a_45200_1800# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X214 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X215 a_17600_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X216 a_5000_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X217 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X218 a_56600_8700# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X219 a_53000_10000# bpa a_52700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X220 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X221 bna en a_8600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X222 ynp znp a_33200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X223 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X224 a_56900_10000# bpa a_56600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X225 avdd bpa a_53000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X226 a_37400_n1600# znp a_37100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X227 a_16100_n1600# bna a_15800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X228 a_23300_10000# zpp a_23000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X229 a_20000_n1600# bna a_19700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X230 a_27200_10000# zpp a_26900_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X231 a_8600_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X232 a_48500_6100# zpp a_48200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X233 a_45200_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X234 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X235 bna_ bnb a_6800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X236 a_200_1800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X237 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X238 a_41600_n3300# bna a_41300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X239 a_45500_n3300# bnb a_45200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X240 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X241 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X242 a_49400_n3300# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X243 a_34100_1800# znp a_33800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X244 a_40400_7400# bpa a_40100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X245 ypm ip a_27800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X246 znp znp a_51800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X247 a_36200_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X248 avss znm a_72800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X249 a_30800_1800# bna a_30500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X250 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X251 a_61400_100# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X252 a_200_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X253 a_43700_n1600# bnb a_43400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X254 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X255 a_47600_n1600# bna a_47300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X256 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X257 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X258 a_53600_100# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X259 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X260 ypm zpp a_29600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X261 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X262 a_30800_6100# zpp a_30500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X263 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X264 a_16100_10000# bpa a_15800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X265 a_20600_100# bna a_20300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X266 a_26600_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X267 a_20000_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X268 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X269 a_23300_7400# zpp a_23000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X270 a_17000_1800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X271 a_56000_1800# znp a_55700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X272 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X273 bnb bnb a_13400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X274 a_45800_100# bnb a_45500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X275 ynp znp a_52400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X276 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X277 ypp zpp a_24800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X278 a_51800_n3300# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X279 a_1700_100# bna a_1400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X280 a_10400_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X281 a_55700_n3300# znp a_55400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X282 a_12800_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X283 avdd zpp a_63800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X284 a_21800_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X285 a_59600_n3300# znp a_59300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X286 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X287 a_8000_1800# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X288 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X289 a_38000_100# znp a_37700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X290 bna_ bnb a_4400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X291 a_17000_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X292 o znm a_71000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X293 a_56000_6100# bpb a_55700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X294 a_1400_1800# bna a_1100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X295 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X296 a_75200_n1600# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X297 a_47300_100# bna a_47000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X298 ynp znp a_53600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X299 a_52700_6100# bpa a_52400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X300 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X301 a_3200_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X302 a_57800_n1600# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X303 bna_ bnb a_14000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X304 a_48500_7400# zpp a_48200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X305 a_20300_n1600# bna a_20000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X306 a_38900_1800# znp a_38600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X307 a_45200_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X308 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X309 a_24200_n1600# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X310 a_8000_6100# bpa a_7700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X311 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X312 a_35600_1800# znp a_35300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X313 a_39500_100# znp a_39200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X314 a_74600_1800# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X315 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X316 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X317 a_32300_1800# znp a_32000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X318 o znm a_71000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X319 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X320 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X321 a_40400_8700# bpa a_40100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X322 a_62000_n3300# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X323 zpm bnb a_65600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X324 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X325 a_69800_n3300# znp a_69500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X326 a_35600_6100# bpa a_35300_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X327 a_200_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X328 a_32300_n3300# znp a_32000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X329 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X330 xp bpa a_32000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X331 a_11000_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X332 a_36200_n3300# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X333 a_14900_n3300# bna a_14600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X334 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X335 a_18800_n3300# bna a_18500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X336 a_18500_1800# bna a_18200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X337 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X338 avss znp a_57200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X339 ypm zpp a_29600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X340 znm bnb a_63800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X341 a_15200_1800# bna a_14900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X342 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X343 a_30800_7400# zpp a_30500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X344 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X345 a_68000_n1600# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X346 a_2000_n3300# bna a_1700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X347 a_60800_100# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X348 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X349 a_54200_1800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X350 a_26600_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X351 bna_ bnb a_5600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X352 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X353 a_30500_n1600# bna a_30200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X354 a_200_n1600# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X355 a_53900_10000# bpa a_53600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X356 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X357 a_9800_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X358 a_34400_n1600# znp a_34100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X359 a_23300_8700# zpp a_23000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X360 a_57800_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X361 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X362 ynm znp a_38000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X363 bna_ bnb a_12800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X364 a_17000_n1600# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X365 bna_ en a_9200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X366 avdd bpa a_20000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X367 a_24200_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X368 a_53000_100# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X369 a_6200_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X370 avdd bpa a_18200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X371 a_1100_n3300# bna a_800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X372 avdd bpa a_57200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X373 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X374 bnb bnb a_3800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X375 zpm bnb a_62000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X376 a_54200_6100# bpa a_53900_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X377 a_8000_n1600# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X378 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X379 a_200_100# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X380 a_17000_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X381 a_56000_7400# bpb a_55700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X382 a_42500_n3300# bna a_42200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X383 bpa_ bpa a_9200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X384 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X385 a_46400_n3300# bnb a_46100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X386 a_52700_7400# bpa a_52400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X387 znp znp a_54200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X388 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X389 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X390 a_48500_8700# zpp a_48200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X391 xn im a_24800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X392 a_29000_n3300# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X393 avss bna a_21200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X394 wn bna a_42800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X395 a_45200_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X396 a_8000_7400# bpa a_7700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X397 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X398 avss znp a_40400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X399 wn bnb a_46400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X400 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X401 avdd zpp a_63800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X402 a_44600_n1600# bnb a_44300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X403 a_2600_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X404 bnb bnb a_13400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X405 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X406 a_48500_n1600# bna a_48200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X407 a_200_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X408 a_30500_10000# zpp a_30200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X409 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X410 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X411 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X412 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X413 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X414 a_38900_100# znp a_38600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X415 a_17000_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X416 a_35600_7400# bpa a_35300_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X417 a_200_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X418 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X419 a_26000_1800# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X420 xp bpa a_32000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X421 a_48200_100# bna a_47900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X422 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X423 a_65000_1800# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X424 a_15200_100# bna a_14900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X425 a_22700_1800# bna a_22400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X426 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X427 a_8000_10000# bpa a_7700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X428 ynp znp a_52400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X429 znm znp a_61400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X430 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X431 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X432 a_56600_n3300# znp a_56300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X433 a_30800_8700# zpp a_30500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X434 a_26000_6100# zpp a_25700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X435 a_72200_n1600# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X436 a_65000_6100# zpp a_64700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X437 a_50900_n1600# znp a_50600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X438 ypp zpp a_22400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X439 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X440 a_54800_n1600# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X441 avdd bpa a_18200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X442 a_58700_n1600# znp a_58400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X443 avdd bpa a_57200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X444 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X445 avdd bpa a_40400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X446 a_21200_n1600# bna a_20900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X447 a_47900_1800# bna a_47600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X448 a_54200_7400# bpa a_53900_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X449 a_44600_10000# zpp a_44300_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X450 a_48500_10000# zpp a_48200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X451 a_44600_1800# bnb a_44300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X452 a_17000_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X453 a_56000_8700# bpb a_55700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X454 a_41300_1800# bna a_41000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X455 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X456 bpa_ bpa a_9200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X457 a_52700_8700# bpa a_52400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X458 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X459 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X460 znm znp a_61400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X461 znm bnb a_62600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X462 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X463 a_8000_8700# bpa a_7700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X464 a_66800_n3300# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X465 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X466 a_44600_6100# zpp a_44300_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X467 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X468 a_33200_n3300# znp a_32900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X469 bna_ bnb a_11600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X470 ynp znp a_53600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X471 a_41300_6100# zpp a_41000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X472 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X473 a_15800_n3300# bna a_15500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X474 a_20900_100# bna a_20600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X475 a_19700_n3300# bna a_19400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X476 a_69800_1800# znp a_69500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X477 ynm znp a_60800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X478 a_63200_100# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X479 xn ip a_27200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X480 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X481 znm bnb a_66200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X482 a_65000_n1600# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X483 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X484 a_30200_100# bna a_29900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X485 a_24200_1800# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X486 bnb bnb a_2600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X487 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X488 a_68900_n1600# znp a_68600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X489 a_63200_1800# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X490 a_35600_8700# bpa a_35300_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X491 a_46100_100# bnb a_45800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X492 a_50900_10000# bpb a_50600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X493 a_6800_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X494 a_31400_n1600# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X495 a_2000_100# bna a_1700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X496 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X497 bna_ bnb a_12800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X498 a_54800_10000# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X499 xp bpa a_32000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X500 a_35300_n1600# znp a_35000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X501 ypm zpp a_58400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X502 a_39200_n1600# znp a_38900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X503 a_14000_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X504 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X505 a_55400_100# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X506 a_21200_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X507 a_17900_n1600# bna a_17600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X508 a_22400_100# bna a_22100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X509 a_69800_6100# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X510 ypm zpp a_27200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X511 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X512 a_24200_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X513 a_5000_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X514 a_63200_6100# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X515 avss znm a_72800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X516 a_47600_100# bna a_47300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X517 bna en a_8600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X518 bna_ bnb a_3200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X519 a_14600_100# bna bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X520 a_26000_7400# zpp a_25700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X521 a_49400_1800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X522 a_65000_7400# zpp a_64700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X523 a_43400_n3300# bnb wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X524 ypp zpp a_22400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X525 a_22100_n3300# bna a_21800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X526 avdd bpa a_18200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X527 a_47300_n3300# bna a_47000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X528 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X529 bna_ bnb a_12800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X530 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X531 a_26000_n3300# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X532 avdd bpa a_57200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X533 a_39800_100# znp a_39500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X534 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X535 znp znp a_51800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X536 a_29900_n3300# bna a_29600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X537 a_54200_8700# bpa a_53900_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X538 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X539 a_41600_n1600# bna a_41300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X540 a_49400_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X541 bpa_ bpa a_9200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X542 a_65000_10000# zpp a_64700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X543 a_45500_n1600# bnb a_45200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X544 bnb bnb a_3800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X545 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X546 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X547 a_49400_n1600# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X548 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X549 a_31400_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X550 ypm ip a_27800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X551 wp bpb a_51800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X552 a_35300_10000# bpa a_35000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X553 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X554 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X555 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X556 avdd bpa a_17600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X557 a_44600_7400# zpp a_44300_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X558 a_41300_7400# zpp a_41000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X559 a_35000_1800# znp a_34700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X560 ynm znp a_60800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X561 a_74000_1800# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X562 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X563 a_31700_1800# znp a_31400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X564 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X565 a_53600_n3300# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X566 avss znp a_70400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X567 a_8900_10000# bpa a_8600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X568 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X569 a_70400_100# znp a_70100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X570 avss znp a_57200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X571 a_40100_n3300# znp a_39800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X572 a_35000_6100# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X573 a_62600_100# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X574 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X575 a_31700_6100# bpa a_31400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X576 a_51800_n1600# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X577 a_69800_7400# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X578 a_55700_n1600# znp a_55400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X579 avdd zpp a_70400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X580 ypm zpp a_27200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X581 a_59600_n1600# znp a_59300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X582 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X583 a_17900_1800# bna a_17600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X584 a_24200_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X585 a_41600_10000# zpp a_41300_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X586 a_63200_7400# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X587 a_56900_1800# znp a_56600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X588 a_45500_10000# zpp a_45200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X589 a_14600_1800# bna bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X590 a_54800_100# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X591 a_49400_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X592 a_53600_1800# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X593 a_26000_8700# zpp a_25700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X594 bnb bnb a_11000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X595 a_28100_10000# zpp a_27800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X596 a_21800_100# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X597 a_65000_8700# zpp a_64700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X598 a_50300_1800# znp a_50000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X599 ypp zpp a_22400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X600 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X601 bna en a_8600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X602 a_47000_100# bna wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X603 a_63800_n3300# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X604 a_5600_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X605 avdd bpa a_17600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X606 bnb bnb a_2600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X607 znm znp a_67400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X608 a_14000_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X609 a_56900_6100# bpa a_56600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X610 bna_ bna a_2000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X611 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X612 a_30200_n3300# bna a_29900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X613 a_56300_100# znp a_56000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X614 a_53600_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X615 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X616 a_49400_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X617 a_23300_100# bna a_23000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X618 wp bpa a_50000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X619 a_12800_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X620 avss bna a_16400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X621 a_39800_1800# znp a_39500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X622 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X623 a_8900_6100# bpa a_8600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X624 a_36500_1800# znp a_36200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X625 a_62000_n1600# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X626 wp bpb a_51800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X627 a_48500_100# bna a_48200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X628 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X629 zpm bnb a_65600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X630 avss znm a_75200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X631 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X632 a_33200_1800# znp a_32900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X633 a_4400_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X634 a_69800_n1600# znp a_69500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X635 a_3800_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X636 a_15500_100# bna a_15200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X637 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X638 a_72200_1800# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X639 a_51800_10000# bpb a_51500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X640 a_44600_8700# zpp a_44300_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X641 bna en a_7400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X642 a_32300_n1600# znp a_32000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X643 a_55700_10000# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X644 a_36200_n1600# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X645 a_11000_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X646 a_41300_8700# zpp a_41000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X647 a_14900_n1600# bna a_14600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X648 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X649 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X650 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X651 a_18800_n1600# bna a_18500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X652 a_39800_6100# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X653 a_36500_6100# bpa a_36200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X654 a_2000_n1600# bna a_1700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X655 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X656 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X657 bna_ bnb a_5600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X658 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X659 a_74000_n3300# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X660 a_9800_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X661 a_19400_1800# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X662 a_35000_7400# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X663 a_40400_n3300# znp a_40100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X664 a_58400_1800# znp a_58100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X665 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X666 a_44300_n3300# bnb a_44000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X667 a_31700_7400# bpa a_31400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X668 a_69800_8700# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X669 ypm zpp a_27200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X670 a_23000_n3300# bna a_22700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X671 a_48200_n3300# bna a_47900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X672 avdd zpp a_70400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X673 a_1100_n1600# bna a_800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X674 ypm ip a_26600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X675 a_22100_1800# bna a_21800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X676 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X677 a_24200_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X678 ynm znp a_60800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X679 a_63200_8700# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X680 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X681 a_62000_100# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X682 a_19400_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X683 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X684 a_42500_n1600# bna a_42200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X685 a_58400_6100# zpp a_58100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X686 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X687 a_46400_n1600# bnb a_46100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X688 o znm a_71000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X689 a_69800_10000# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X690 xn im a_24800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X691 a_22100_6100# zpp a_21800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X692 xp bpa a_32000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X693 a_29000_n1600# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X694 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X695 avdd bpa a_17600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X696 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X697 a_36200_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X698 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X699 a_56900_7400# bpa a_56600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X700 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X701 a_18800_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X702 a_53600_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X703 zpm bnb a_63200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X704 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X705 a_49400_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X706 a_44000_1800# bnb a_43700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X707 wp bpa a_50000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X708 a_30500_100# bna a_30200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X709 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X710 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X711 a_50600_n3300# znp a_50300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X712 avss znp a_40400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X713 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X714 a_8900_7400# bpa a_8600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X715 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X716 wp bpb a_51800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X717 znp znp a_54200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X718 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X719 a_58400_n3300# znp a_58100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X720 a_55700_100# znp a_55400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X721 a_37100_n3300# znp a_36800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X722 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X723 a_22700_100# bna a_22400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X724 bpa_ bpa a_800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X725 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X726 a_44000_6100# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X727 a_39800_7400# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X728 ynp znp a_52400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X729 a_47900_100# bna a_47600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X730 avdd bpa a_40400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X731 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X732 a_3800_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X733 a_36500_7400# bpa a_36200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X734 a_56600_n1600# znp a_56300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X735 a_14900_100# bna a_14600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X736 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X737 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X738 a_57200_100# znp a_56900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X739 ypm ip a_26600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X740 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X741 zpm bnb a_65600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X742 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X743 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X744 a_23600_1800# bna a_23300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X745 a_24200_100# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X746 ypp zpp a_24800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X747 a_40100_100# znp a_39800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X748 a_62600_1800# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X749 a_35000_8700# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X750 a_20300_1800# bna a_20000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X751 a_29000_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X752 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X753 a_500_1800# bna a_200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X754 a_31700_8700# bpa a_31400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X755 avdd zpp a_70400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X756 a_49400_100# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X757 bnb bnb a_5000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X758 a_60800_n3300# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X759 a_16400_100# bna a_16100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X760 a_26900_6100# zpp a_26600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X761 zpm bnb a_64400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X762 a_68600_n3300# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X763 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X764 a_23600_6100# zpp a_23300_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X765 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X766 a_19400_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X767 avdd bpa a_20000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X768 a_58400_7400# zpp a_58100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X769 bnb bnb a_13400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X770 a_500_6100# bpa a_200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X771 a_17600_n3300# bna a_17300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X772 a_48800_1800# bna a_48500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X773 a_22100_7400# zpp a_21800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X774 znm bnb a_62600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X775 a_45500_1800# bnb a_45200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X776 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X777 avdd bpa a_17600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X778 a_56900_8700# bpa a_56600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X779 a_66800_n1600# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X780 a_42200_1800# bna a_41900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X781 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X782 bna_ bnb a_4400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X783 a_53600_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X784 a_52700_10000# bpa a_52400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X785 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X786 a_8600_n3300# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X787 a_33200_n1600# znp a_32900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X788 a_56600_10000# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X789 bna_ bnb a_11600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X790 avss znp a_70400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X791 wp bpa a_50000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X792 a_15800_n1600# bna a_15500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X793 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X794 a_19700_n1600# bna a_19400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X795 a_8900_8700# bpa a_8600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X796 a_48800_6100# zpp a_48500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X797 a_45500_6100# zpp a_45200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X798 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X799 bnb bnb a_2600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X800 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X801 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X802 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X803 a_71000_n3300# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X804 znm bnb a_62600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X805 a_6800_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X806 o znm a_74600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X807 a_28400_1800# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X808 a_72200_100# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X809 a_44000_7400# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X810 a_41300_n3300# bna a_41000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X811 a_67400_1800# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X812 a_39800_8700# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X813 a_45200_n3300# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X814 avdd bpa a_40400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X815 xn bna a_23600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X816 ynp znp a_54800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X817 a_36500_8700# bpa a_36200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X818 avss bna a_30800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X819 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X820 a_27800_n3300# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X821 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X822 a_22100_100# bna a_21800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X823 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X824 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X825 avss znm a_72800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X826 a_64400_100# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X827 a_31400_100# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X828 a_28400_6100# zpp a_28100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X829 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X830 a_43400_n1600# bnb wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X831 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X832 a_22100_n1600# bna a_21800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X833 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X834 a_47300_n1600# bna a_47000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X835 a_26000_n1600# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X836 a_56600_100# znp a_56300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X837 avdd zpp a_30800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X838 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X839 a_29900_n1600# bna a_29600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X840 a_23600_100# bna a_23300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X841 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X842 a_26900_7400# zpp a_26600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X843 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X844 a_15800_10000# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X845 a_23600_7400# zpp a_23300_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X846 avdd bpa a_19400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X847 a_19400_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X848 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X849 avdd bpa a_20000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X850 a_14000_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X851 a_58400_8700# zpp a_58100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X852 a_48800_100# bna a_48500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X853 a_500_7400# bpa a_200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X854 a_53000_1800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X855 bna_ bnb a_4400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X856 bna_ bnb a_10400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X857 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X858 a_15800_100# bna a_15500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X859 ynp znp a_51200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X860 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X861 a_22100_8700# zpp a_21800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X862 a_55400_n3300# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X863 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X864 a_34100_n3300# znp a_33800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X865 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X866 a_59300_n3300# znp a_59000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X867 a_38000_n3300# znp a_37700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X868 a_5000_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X869 a_1700_1800# bna a_1400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X870 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X871 a_53000_6100# bpa a_52700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X872 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X873 a_6200_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X874 a_17300_100# bna a_17000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X875 a_48800_7400# zpp a_48500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X876 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X877 a_53600_n1600# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X878 avss znp a_57200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X879 a_45500_7400# zpp a_45200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X880 avss znp a_35600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X881 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X882 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X883 a_40100_n1600# znp a_39800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X884 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X885 a_22100_10000# zpp a_21800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X886 o znm a_74600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X887 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X888 a_32600_1800# znp a_32300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X889 a_26000_10000# zpp a_25700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X890 a_71600_1800# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X891 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X892 a_44000_8700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X893 ypm zpp a_29600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X894 avdd bpa a_40400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X895 znm znp a_61400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X896 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X897 a_65600_n3300# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X898 avdd bpa a_35600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X899 a_71600_100# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X900 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X901 a_69500_n3300# znp a_69200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X902 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X903 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X904 a_28400_7400# zpp a_28100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X905 bna_ bnb a_10400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X906 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X907 a_14600_n3300# bna bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X908 a_18800_1800# bna a_18500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X909 a_18500_n3300# bna a_18200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X910 a_57800_1800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X911 a_15500_1800# bna a_15200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X912 avdd zpp a_30800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X913 a_63800_100# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X914 a_63800_n1600# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X915 znp znp a_54200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X916 a_26900_8700# zpp a_26600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X917 a_12200_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X918 a_30800_100# bna a_30500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X919 znm znp a_67400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X920 a_1700_n3300# bna a_1400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X921 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X922 a_51200_1800# znp a_50900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X923 a_23600_8700# zpp a_23300_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X924 a_5600_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X925 a_30200_n1600# bna a_29900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X926 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X927 a_53600_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X928 bna_ en a_9200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X929 avdd bpa a_20000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X930 a_9800_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X931 avdd bpa a_57200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X932 a_500_8700# bpa a_200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X933 a_12800_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X934 a_56000_100# znp a_55700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X935 avss bna a_16400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X936 bnb bnb a_6200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X937 a_18800_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X938 a_40100_10000# bpa a_39800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X939 a_23000_100# bna a_22700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X940 a_57800_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X941 a_3200_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X942 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X943 a_800_n3300# bna a_500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X944 znm bnb a_65000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X945 wp bpa a_54200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X946 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X947 a_3800_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X948 a_32300_100# znp a_32000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X949 znp bpb a_50900_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X950 avss znm a_71600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X951 bna en a_7400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X952 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X953 bnb bnb a_3800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X954 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X955 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X956 a_37400_1800# znp a_37100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X957 a_53000_7400# bpa a_52700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X958 a_42200_n3300# bna a_41900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X959 avss znp a_57200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X960 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X961 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X962 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X963 a_48800_8700# zpp a_48500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X964 a_20900_n3300# bna a_20600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X965 ypp im a_24200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X966 a_24800_n3300# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X967 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X968 a_45500_8700# zpp a_45200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X969 xn ip a_28400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X970 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X971 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X972 a_74000_n1600# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X973 a_49700_100# znp a_49400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X974 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X975 a_5600_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X976 a_40400_n1600# znp a_40100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X977 avss bna a_16400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X978 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X979 a_63800_10000# zpp a_63500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X980 a_44300_n1600# bnb a_44000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X981 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X982 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X983 a_48200_n1600# bna a_47900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X984 a_23000_n1600# bna a_22700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X985 ypm ip a_26600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X986 a_30200_10000# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X987 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X988 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X989 avdd bpa a_35600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X990 a_59300_1800# znp a_59000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X991 avdd bpa a_16400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X992 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X993 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X994 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X995 a_28400_8700# zpp a_28100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X996 a_18200_100# bna a_17900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X997 a_23000_1800# bna a_22700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X998 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X999 a_62000_1800# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1000 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1001 a_7700_10000# bpa a_7400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1002 a_52400_n3300# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1003 avdd zpp a_30800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1004 avss bna a_30800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1005 a_56300_n3300# znp a_56000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1006 a_71000_100# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1007 a_35000_n3300# znp a_34700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1008 a_38900_n3300# znp a_38600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1009 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1010 a_23000_6100# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1011 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1012 a_18800_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1013 a_50600_n1600# znp a_50300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1014 a_57800_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1015 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1016 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1017 znp znp a_54200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1018 a_58400_n1600# znp a_58100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1019 wp bpa a_54200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1020 o znm a_72200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1021 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1022 a_40400_10000# bpa a_40100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1023 a_37100_n1600# znp a_36800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1024 zpp bnb a_44600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1025 znp bpb a_50900_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1026 a_44300_10000# zpp a_44000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1027 a_23000_10000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1028 a_48200_10000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1029 a_41600_1800# bna a_41300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1030 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1031 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1032 a_26900_10000# zpp a_26600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1033 a_53000_8700# bpa a_52700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1034 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1035 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1036 zpm bnb a_64400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1037 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1038 a_31700_100# znp a_31400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1039 a_62600_n3300# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1040 avdd zpp a_44600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1041 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1042 znm bnb a_66200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1043 a_56900_100# znp a_56600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1044 a_41600_6100# zpp a_41300_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1045 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1046 avss bna a_48800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1047 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1048 a_11600_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1049 xn bna a_23600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1050 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1051 a_70100_1800# znp a_69800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1052 a_15500_n3300# bna a_15200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1053 a_66200_100# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1054 a_27800_1800# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1055 a_19400_n3300# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1056 a_66800_1800# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1057 a_60800_n1600# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1058 a_33200_100# znp a_32900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1059 ypp im a_24200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1060 zpm bnb a_63200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1061 avdd bpa a_35600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1062 zpm bnb a_64400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1063 avss bna a_48800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1064 a_21200_1800# bna a_20900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1065 a_68600_n1600# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1066 a_2600_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1067 a_5000_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1068 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1069 a_60200_1800# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1070 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1071 a_16100_100# bna a_15800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1072 a_50600_10000# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1073 bnb bnb a_6200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1074 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1075 a_58400_100# znp a_58100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1076 wp bpa a_54200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1077 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1078 a_58400_10000# zpp a_58100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1079 bnb bnb a_13400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1080 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1081 a_25400_100# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1082 a_70100_6100# zpp a_69800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1083 xp bpa a_36800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1084 a_17600_n1600# bna a_17300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1085 a_27800_6100# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1086 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1087 a_24500_6100# zpp a_24200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1088 a_63500_6100# zpp a_63200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1089 a_21200_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1090 bna_ bnb a_4400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1091 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1092 bnb bnb a_6200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1093 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1094 a_72800_n3300# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1095 a_17600_100# bna a_17300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1096 a_8600_n1600# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1097 a_49700_1800# znp a_49400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1098 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X1099 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1100 a_23000_7400# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1101 a_46400_1800# bnb a_46100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1102 a_18800_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1103 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1104 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1105 a_57800_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1106 a_21800_n3300# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1107 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1108 wp bpa a_54200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1109 ypp im a_25400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1110 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1111 a_29600_n3300# bna a_29300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1112 znp bpb a_50900_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1113 a_71000_n1600# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1114 o znm a_74600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1115 a_49700_6100# bpa a_49400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1116 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1117 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1118 a_41300_n1600# bna a_41000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1119 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1120 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1121 a_64700_10000# zpp a_64400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1122 a_45200_n1600# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1123 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1124 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1125 xn bna a_23600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1126 avss znm a_71600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1127 a_27800_n1600# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1128 a_29300_1800# bna a_29000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1129 avdd zpp a_44600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1130 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1131 ynm znp a_68000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1132 a_17600_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1133 a_41600_7400# zpp a_41300_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1134 znm bnb a_63800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1135 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1136 a_32000_1800# znp a_31700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1137 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X1138 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1139 avss bna a_30800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1140 a_71000_1800# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1141 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1142 a_73400_100# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1143 znp znp a_53000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1144 a_8600_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1145 a_32000_n3300# znp a_31700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1146 a_40400_100# znp a_40100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1147 a_57200_n3300# znp a_56900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1148 a_29300_6100# zpp a_29000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1149 avss znp a_35600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1150 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1151 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1152 a_39800_n3300# znp a_39500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1153 a_65600_100# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1154 a_32000_6100# bpa a_31700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1155 a_70100_7400# zpp a_69800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1156 a_32600_100# znp a_32300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1157 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1158 a_27800_7400# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1159 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1160 ynp znp a_51200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1161 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1162 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1163 a_55400_n1600# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1164 a_24500_7400# zpp a_24200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1165 a_34100_n1600# znp a_33800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1166 a_63500_7400# zpp a_63200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1167 a_59300_n1600# znp a_59000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1168 a_14900_1800# bna a_14600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1169 a_21200_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1170 a_41300_10000# zpp a_41000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1171 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1172 a_38000_n1600# znp a_37700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1173 a_57800_100# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1174 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1175 ynp znp a_53600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1176 a_45200_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1177 a_11600_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1178 a_24800_100# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1179 avdd zpp a_23600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1180 a_50600_1800# znp a_50300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1181 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1182 a_23000_8700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1183 a_27800_10000# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1184 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1185 a_50000_100# znp a_49700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1186 bna_ bnb a_5600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1187 bna_ bnb a_5600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1188 a_17000_100# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1189 zpm bnb a_63200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1190 a_2600_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1191 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1192 a_59300_100# znp a_59000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1193 a_53900_6100# bpa a_53600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1194 a_67400_n3300# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1195 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1196 a_46100_n3300# bnb a_45800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1197 a_49700_7400# bpa a_49400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1198 xn im a_26000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1199 a_50600_6100# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1200 a_50000_n3300# znp a_49700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1201 a_40100_1800# znp a_39800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1202 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1203 bnb bnb a_12200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1204 a_16400_n3300# bna a_16100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1205 a_36800_1800# znp a_36500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1206 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1207 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1208 ynp znp a_33200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1209 znm znp a_61400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1210 a_7400_100# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1211 a_18500_100# bna a_18200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1212 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1213 a_65600_n1600# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1214 o znm a_72200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1215 avdd zpp a_44600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1216 a_30200_1800# bna a_29900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1217 bna_ bnb a_3200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1218 a_69500_n1600# znp a_69200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1219 a_51500_10000# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1220 a_41600_8700# zpp a_41300_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1221 a_7400_n3300# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1222 znp bpb a_55100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1223 bna_ bnb a_10400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1224 a_40100_6100# bpa a_39800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1225 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1226 a_14600_n1600# bna bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1227 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1228 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1229 a_18500_n1600# bna a_18200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1230 a_36800_6100# bpa a_36500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1231 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1232 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1233 a_1700_n1600# bna a_1400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1234 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1235 a_29300_7400# zpp a_29000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1236 a_30200_6100# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1237 a_5600_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1238 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1239 a_19700_1800# bna a_19400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1240 o znm a_73400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1241 bna_ en a_9200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1242 a_58700_1800# znp a_58400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1243 a_16400_1800# bna a_16100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1244 a_72800_100# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1245 a_32000_7400# bpa a_31700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1246 a_70100_8700# zpp a_69800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1247 a_55400_1800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1248 a_27800_8700# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1249 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1250 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1251 a_24500_8700# zpp a_24200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1252 a_22700_n3300# bna a_22400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1253 a_800_n1600# bna a_500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1254 a_26600_n3300# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1255 a_63500_8700# zpp a_63200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1256 a_21200_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1257 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1258 avss znm a_71600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1259 a_65000_100# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1260 a_7400_1800# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1261 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1262 avdd bpa a_19400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1263 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1264 a_32000_100# znp a_31700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1265 ypm zpp a_58400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1266 a_16400_6100# bpa a_16100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1267 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1268 a_42200_n1600# bna a_41900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1269 avss znm a_74000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1270 znp bpb a_55100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1271 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1272 a_20900_n1600# bna a_20600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1273 a_41300_100# bna a_41000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1274 a_24800_n1600# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1275 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1276 xn ip a_28400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1277 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1278 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1279 ynm znp a_38000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1280 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1281 a_53900_7400# bpa a_53600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1282 znm bnb a_66200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1283 a_7400_6100# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1284 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1285 avdd bpa a_18200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1286 a_49700_8700# bpa a_49400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1287 a_50600_7400# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1288 ynp znp a_33200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1289 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1290 a_41000_1800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1291 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1292 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1293 a_50300_n3300# znp a_50000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1294 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1295 a_58700_100# znp a_58400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1296 bpa_ bpa a_9200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1297 a_54200_n3300# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1298 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1299 a_32900_n3300# znp a_32600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1300 ypp im a_25400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1301 a_36800_n3300# znp a_36500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1302 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1303 a_800_10000# bpa a_500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1304 a_40100_7400# bpa a_39800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1305 a_41000_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1306 a_6800_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1307 a_36800_7400# bpa a_36500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1308 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1309 a_52400_n1600# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1310 a_17900_100# bna a_17600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1311 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1312 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1313 a_56300_n1600# znp a_56000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1314 avss bna a_30800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1315 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1316 a_29300_8700# zpp a_29000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1317 a_35000_n1600# znp a_34700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1318 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1319 xn bna a_23600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1320 a_30200_7400# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1321 a_38900_n1600# znp a_38600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1322 a_27200_100# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1323 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1324 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1325 znm bnb a_62600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1326 avdd bpa a_20600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1327 a_20600_1800# bna a_20300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1328 a_24800_10000# zpp a_24500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1329 a_800_1800# bna a_500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1330 a_32000_8700# bpa a_31700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1331 avdd zpp a_28400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1332 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1333 bna_ en a_8000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1334 a_19400_100# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1335 znm znp a_60200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1336 avdd zpp a_23600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1337 a_64400_n3300# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1338 wn bna a_42800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1339 ynm znp a_68000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1340 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1341 avdd bpa a_19400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1342 a_20600_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1343 a_47000_n3300# bna wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1344 ypm zpp a_58400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1345 a_800_6100# bpa a_500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1346 a_16400_7400# bpa a_16100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1347 znp bpb a_55100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1348 avss bna a_48800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1349 a_13400_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1350 a_500_100# bna a_200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1351 a_17300_n3300# bna a_17000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1352 a_45800_1800# bnb a_45500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1353 a_42500_1800# bna a_42200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1354 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1355 a_62600_n1600# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1356 a_53900_8700# bpa a_53600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1357 znm bnb a_66200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1358 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1359 a_4400_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1360 a_7400_7400# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1361 o znm a_73400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1362 a_50600_8700# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1363 avss bna a_48800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1364 bna_ en a_8000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1365 a_52400_10000# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1366 avdd zpp a_30800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1367 wp bpb a_56000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1368 a_11600_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1369 avss znp a_40400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1370 avdd zpp a_48800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1371 a_35000_10000# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1372 a_15500_n1600# bna a_15200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1373 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1374 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1375 a_19400_n1600# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1376 a_45800_6100# zpp a_45500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1377 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1378 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1379 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1380 zpm bnb a_65600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1381 a_2600_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1382 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1383 a_32900_100# znp a_32600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1384 avss znp a_70400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1385 bnb bnb a_6200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1386 xn ip a_28400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1387 a_74600_n3300# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1388 a_75200_100# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1389 znm znp a_67400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1390 a_40100_8700# bpa a_39800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1391 a_42200_100# bna a_41900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1392 a_25400_1800# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1393 a_41000_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1394 a_58100_100# znp a_57800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1395 a_64400_1800# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1396 a_36800_8700# bpa a_36500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1397 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1398 a_23600_n3300# bna a_23300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1399 xn im a_24800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1400 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1401 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1402 xn ip a_27200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1403 a_67400_100# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1404 a_30200_8700# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1405 a_72800_n1600# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1406 a_34400_100# znp a_34100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1407 avdd zpp a_28400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1408 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X1409 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1410 a_25400_6100# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1411 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1412 a_64400_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1413 a_21800_n1600# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1414 a_59600_100# znp a_59300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1415 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1416 ypp im a_25400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1417 a_26600_100# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1418 avdd zpp a_48800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1419 a_29600_n1600# bna a_29300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1420 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1421 avdd zpp a_23600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1422 a_47300_1800# bna a_47000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1423 avdd bpa a_19400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1424 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1425 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1426 a_20600_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1427 a_19400_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1428 ypm zpp a_58400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1429 a_16400_8700# bpa a_16100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1430 a_800_7400# bpa a_500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1431 bna en a_7400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1432 a_11000_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1433 znp bpb a_55100_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1434 a_18800_100# bna a_18500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1435 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1436 a_51200_n3300# znp a_50900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1437 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1438 a_33800_n3300# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1439 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1440 a_7400_8700# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1441 a_37700_n3300# znp a_37400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1442 a_2000_1800# bna a_1700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1443 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1444 a_9200_100# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1445 avdd zpp a_48800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1446 a_45800_7400# zpp a_45500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1447 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1448 znp znp a_53000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1449 a_69200_1800# znp a_68900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1450 a_32000_n1600# znp a_31700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1451 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X1452 a_57200_n1600# znp a_56900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1453 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1454 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1455 avss znp a_35600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1456 avss znm a_72800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1457 a_32900_1800# znp a_32600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1458 a_39800_n1600# znp a_39500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1459 avss znm a_71600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1460 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1461 a_21800_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1462 a_25700_10000# zpp a_25400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1463 a_41000_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1464 a_29600_10000# zpp a_29300_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1465 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1466 a_61400_n3300# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1467 a_74600_100# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1468 znm bnb a_65000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1469 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1470 a_44000_n3300# bnb a_43700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1471 a_41600_100# bna a_41300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1472 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1473 avdd zpp a_28400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1474 a_69200_n3300# znp a_68900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1475 a_47900_n3300# bna a_47600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1476 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1477 a_25400_7400# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1478 bpb bna a_18800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1479 a_10400_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1480 a_58100_1800# znp a_57800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1481 a_64400_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1482 bna_ bnb a_14000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1483 a_15800_1800# bna a_15500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1484 a_66800_100# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1485 a_18200_n3300# bna a_17900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1486 a_54800_1800# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1487 bnb bnb a_12200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1488 a_33800_100# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1489 zpm bnb a_63200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1490 ynp znp a_51200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1491 avdd zpp a_23600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1492 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1493 a_67400_n1600# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1494 a_1400_n3300# bna a_1100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1495 a_20600_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1496 a_46100_n1600# bnb a_45800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1497 bnb bnb a_5000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1498 bnb bnb a_9800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1499 a_800_8700# bpa a_500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1500 avdd bpa a_53000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1501 a_50000_n1600# znp a_49700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1502 a_9200_n3300# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1503 a_59000_100# znp a_58700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1504 a_6800_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1505 avdd bpa a_18800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1506 a_32000_10000# bpa a_31700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1507 bnb bnb a_12200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1508 a_57200_10000# bpa a_56900_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1509 a_26000_100# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1510 a_58100_6100# zpp a_57800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1511 avdd bpa a_35600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1512 a_16400_n1600# bna a_16100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1513 bna_ bnb a_3200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1514 a_15800_6100# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1515 ynm znp a_68000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1516 a_39800_10000# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1517 a_54800_6100# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1518 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1519 a_500_n3300# bna a_200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1520 a_35300_100# znp a_35000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1521 a_51500_6100# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1522 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1523 bna_ bnb a_3200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1524 bna_ bnb a_6800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1525 a_71600_n3300# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1526 a_7400_n1600# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1527 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1528 avss znm a_75200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1529 a_37700_1800# znp a_37400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1530 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X1531 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1532 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1533 avdd zpp a_48800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1534 a_34400_1800# znp a_34100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1535 a_58100_n3300# znp a_57800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1536 xn ip a_27200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1537 a_73400_1800# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1538 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1539 a_45800_8700# zpp a_45500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1540 a_20600_n3300# bna a_20300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1541 ypp im a_24200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1542 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1543 a_28400_n3300# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1544 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1545 o znm a_73400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1546 a_8600_100# en bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1547 a_19700_100# bna a_19400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1548 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1549 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X1550 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1551 a_63500_10000# zpp a_63200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1552 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1553 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1554 a_22700_n1600# bna a_22400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1555 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1556 ypp zpp a_45800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1557 a_26600_n1600# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1558 a_50000_10000# bpa a_49700_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1559 a_59600_1800# znp a_59300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1560 a_17300_1800# bna a_17000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1561 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1562 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1563 a_800_100# bna a_500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1564 a_56300_1800# znp a_56000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1565 a_16400_10000# bpa a_16100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1566 avdd zpp a_28400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1567 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1568 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1569 a_25400_8700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1570 a_64400_8700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1571 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1572 a_74000_100# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1573 a_7400_10000# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1574 bna_ en a_8000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1575 a_30800_n3300# bna a_30500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1576 a_41000_100# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1577 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1578 avdd bpa a_17000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1579 a_34700_n3300# znp a_34400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1580 wp bpb a_56000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1581 a_38600_n3300# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1582 a_50300_100# znp a_50000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1583 avdd bpa a_18800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1584 a_58100_7400# zpp a_57800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1585 a_15800_7400# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1586 a_50300_n1600# znp a_50000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1587 a_39200_1800# znp a_38900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1588 a_54800_7400# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1589 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1590 avss znm a_75200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1591 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1592 a_54200_n1600# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1593 avdd bpa a_8000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1594 a_32900_n1600# znp a_32600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1595 a_51500_7400# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1596 a_42500_100# bna a_42200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1597 a_36800_n1600# znp a_36500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1598 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1599 a_41900_1800# bna a_41600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1600 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1601 ypp zpp a_22400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1602 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1603 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1604 a_26600_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1605 znm znp a_67400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1606 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1607 a_34700_100# znp a_34400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1608 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1609 zpm bnb a_62000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1610 a_41000_n3300# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1611 a_66200_n3300# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1612 ynm znp a_59600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1613 ypp zpp a_41600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1614 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1615 zpp bnb a_44600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1616 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1617 ypm ip a_26600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1618 a_48800_n3300# bna a_48500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1619 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X1620 a_69200_100# znp a_68900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1621 ypm ip a_27800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1622 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1623 bnb bnb a_11000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1624 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1625 ynm znp a_66800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1626 a_15200_n3300# bna a_14900_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1627 a_36200_100# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1628 a_24800_1800# im ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1629 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1630 a_63800_1800# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1631 znm znp a_60200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1632 avss bna a_21200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1633 a_8000_100# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1634 znm znp a_60200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1635 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1636 a_64400_n1600# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1637 bpb bna a_18800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1638 wn bna a_42800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1639 ynm znp a_68000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1640 bna_ bna a_2000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1641 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1642 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1643 wp bpa a_50000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1644 a_47000_n1600# bna wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1645 a_6200_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1646 a_54200_10000# bpa a_53900_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1647 a_28400_100# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1648 a_28100_6100# zpp a_27800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1649 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1650 a_13400_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1651 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1652 a_36800_10000# bpa a_36500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1653 a_17300_n1600# bna a_17000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1654 a_24800_6100# zpp a_24500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1655 a_63800_6100# zpp a_63500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1656 avdd bpa a_21200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1657 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1658 bna_ en a_9200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1659 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1660 avdd bpa a_17000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1661 a_4400_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1662 a_50000_1800# znp a_49700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1663 wp bpb a_56000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1664 o znm a_72200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1665 bna_ en a_8000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1666 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1667 wn bnb a_46400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1668 avdd bpa a_18800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1669 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1670 ynp znp a_54800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1671 a_58100_8700# zpp a_57800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1672 a_43400_1800# bnb wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1673 a_15800_8700# bpa bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1674 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1675 a_59000_n3300# znp a_58700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1676 a_54800_8700# bpb wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1677 avss bna a_21200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1678 bpa_ enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1679 avdd bpa a_8000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1680 a_51500_8700# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1681 a_25400_n3300# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1682 a_29300_n3300# bna a_29000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1683 avss znp a_70400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1684 a_50000_6100# bpa a_49700_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1685 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1686 a_74600_n1600# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1687 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1688 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1689 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1690 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1691 o znm a_74600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1692 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1693 a_64400_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1694 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1695 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1696 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1697 a_23600_n1600# bna a_23300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1698 a_41900_100# bna a_41600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1699 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1700 xn ip a_27200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1701 a_29600_1800# bna a_29300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1702 a_68600_1800# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1703 xn im a_26000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1704 a_51200_100# znp a_50900_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1705 ypp zpp a_41600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1706 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1707 ynm znp a_66800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1708 znm bnb a_65000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1709 avdd bpa a_17000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1710 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1711 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X1712 a_34100_100# znp a_33800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1713 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1714 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1715 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1716 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1717 a_43400_100# bnb wn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1718 avdd bpa a_8000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1719 a_29600_6100# zpp a_29300_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1720 a_31700_n3300# znp a_31400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1721 a_10400_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1722 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1723 avdd zpp a_26000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1724 a_35600_n3300# znp a_35300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1725 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1726 ypm zpp a_65000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1727 a_39500_n3300# znp a_39200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1728 a_68600_100# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1729 a_35600_100# znp a_35300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1730 a_28100_7400# zpp a_27800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1731 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1732 a_24800_7400# zpp a_24500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1733 avdd zpp a_70400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1734 a_51200_n1600# znp a_50900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1735 a_48200_1800# bna a_47900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1736 a_63800_7400# zpp a_63500_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1737 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1738 avdd bpa a_21200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1739 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1740 a_33800_n1600# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1741 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1742 avdd bpa a_17000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1743 bna_ bnb a_11600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1744 wp bpb a_56000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1745 a_37700_n1600# znp a_37400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1746 a_27800_100# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1747 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1748 a_50900_1800# znp a_50600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1749 a_23600_10000# zpp a_23300_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1750 ypm zpp a_27200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1751 bna en a_8600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1752 a_48200_6100# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1753 avdd bpa a_8000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1754 a_20000_100# bna a_19700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1755 bnb bnb a_2600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1756 a_63200_n3300# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1757 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1758 a_50000_7400# bpa a_49700_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1759 a_41900_n3300# bna a_41600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1760 a_29300_100# bna a_29000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1761 a_50900_6100# bpb a_50600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1762 a_45800_n3300# bnb a_45500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1763 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1764 a_49700_n3300# znp a_49400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1765 a_37100_1800# znp a_36800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1766 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1767 a_12200_n3300# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1768 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1769 a_1100_100# bna a_800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1770 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1771 a_33800_1800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1772 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1773 a_72800_1800# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1774 a_61400_n1600# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1775 a_30500_1800# bna a_30200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1776 znm bnb a_65000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1777 ypp zpp a_41600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1778 a_44000_n1600# bnb a_43700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1779 a_3200_n3300# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1780 a_69200_n1600# znp a_68900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1781 znp bpb a_50900_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1782 a_47900_n1600# bna a_47600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1783 a_10400_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1784 xp bpa a_36800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1785 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1786 bna_ bnb a_14000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1787 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1788 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1789 a_18200_n1600# bna a_17900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1790 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1791 a_50600_100# znp a_50300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1792 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1793 a_29600_7400# zpp a_29300_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1794 a_30500_6100# zpp a_30200_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1795 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1796 a_1400_n1600# bna a_1100_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1797 a_20000_1800# bna a_19700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1798 avdd zpp a_26000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1799 bnb bnb a_5000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1800 ypm zpp a_65000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1801 a_59000_1800# znp a_58700_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1802 a_73400_n3300# znm avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1803 avss bna a_16400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1804 a_9200_n1600# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1805 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1806 a_55700_1800# znp a_55400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1807 a_28100_8700# zpp a_27800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1808 znp znp a_51800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1809 a_13400_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1810 a_56000_n3300# znp a_55700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1811 a_42800_100# bna a_42500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1812 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1813 a_52400_1800# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1814 a_24800_8700# zpp a_24500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1815 ynm znp a_59600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1816 a_63800_8700# zpp a_63500_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1817 a_22400_n3300# bna a_22100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1818 avdd bpa a_21200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1819 a_500_n1600# bna a_200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1820 xn im a_26000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1821 znm bpb zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1822 a_68000_100# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1823 bna en a_7400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1824 a_20000_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1825 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1826 a_71600_n1600# znm o avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1827 a_35000_100# znp a_34700_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1828 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1829 a_4400_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1830 avss znm a_75200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1831 avdd bpa a_16400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1832 a_55700_6100# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1833 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1834 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1835 a_58100_n1600# znp a_57800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1836 a_44300_100# bnb a_44000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1837 a_52400_6100# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1838 ypm zpp a_65000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1839 a_20600_n1600# bna a_20300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1840 bnb bnb a_11000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1841 a_48200_7400# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1842 a_44000_10000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1843 ypp im a_24200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1844 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1845 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1846 a_28400_n1600# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1847 a_38600_1800# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1848 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1849 a_69500_100# znp a_69200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1850 a_7700_6100# bpa a_7400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1851 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1852 a_50000_8700# bpa a_49700_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1853 a_35300_1800# znp a_35000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1854 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1855 a_50900_7400# bpb a_50600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1856 a_36500_100# znp a_36200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1857 avss znm a_74000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1858 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1859 ypp zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1860 a_18200_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1861 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1862 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1863 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1864 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1865 a_70100_n3300# znp a_69800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1866 xn ip a_28400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1867 a_9200_10000# bpa a_8900_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1868 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1869 a_32600_n3300# znp a_32300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1870 a_36500_n3300# znp a_36200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1871 a_35300_6100# bpa a_35000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1872 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1873 bpb bna a_18800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1874 a_500_10000# bpa a_200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1875 a_9800_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1876 xp bpa a_36800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1877 a_18200_1800# bna a_17900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1878 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1879 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1880 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1881 a_57200_1800# znp a_56900_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1882 a_29600_8700# zpp a_29300_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1883 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1884 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1885 a_30800_n1600# bna a_30500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1886 a_30500_7400# zpp a_30200_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1887 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1888 bnb bnb a_9800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1889 avdd zpp a_26000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1890 a_34700_n1600# znp a_34400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1891 a_20900_1800# bna a_20600_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1892 a_58100_10000# zpp a_57800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1893 a_38600_n1600# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1894 ypm zpp a_65000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1895 a_1100_1800# bna a_800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1896 a_20600_10000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1897 a_24500_10000# zpp a_24200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1898 a_9200_1800# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1899 a_28400_10000# zpp a_28100_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1900 a_18200_6100# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1901 a_57200_6100# bpa a_56900_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1902 a_60200_n3300# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1903 a_20000_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1904 avdd bpa a_20600_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1905 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1906 a_42800_n3300# bna a_42500_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1907 bpa_ bpa a_800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1908 avdd bpa a_16400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1909 wn bnb a_46400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1910 a_55700_7400# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1911 a_9200_6100# bpa a_8900_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1912 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1913 a_52400_7400# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1914 a_46100_1800# bnb a_45800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1915 ynp znp a_51200_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1916 a_48200_8700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1917 a_42800_1800# bna a_42500_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1918 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1919 zpm bnb a_62000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1920 a_7700_7400# bpa a_7400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1921 a_41000_n1600# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1922 a_66200_n1600# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1923 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X1924 a_50900_8700# bpb a_50600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1925 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1926 zpp bnb a_44600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1927 a_43700_100# bnb a_43400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1928 a_48800_n1600# bna a_48500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1929 a_30800_10000# zpp a_30500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1930 bnb bnb a_11000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1931 bna_ bnb a_10400_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1932 ypp zpp a_45800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1933 xp ip ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1934 a_15200_n1600# bna a_14900_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1935 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1936 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1937 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1938 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1939 a_68900_100# znp a_68600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1940 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1941 avss znp a_35600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1942 bna_ bna a_2000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1943 a_29000_1800# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1944 a_35300_7400# bpa a_35000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1945 a_70400_n3300# znp a_70100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1946 a_6200_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1947 a_68000_1800# znp znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1948 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1949 ypp im a_25400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1950 avss znm a_74000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1951 a_45200_100# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1952 a_53000_n3300# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1953 zpm bnb a_64400_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1954 xp bpa a_36800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1955 a_12200_100# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1956 a_22400_1800# bna a_22100_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1957 avdd en zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1958 a_56900_n3300# znp a_56600_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1959 ypm ip a_27800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1960 a_61400_1800# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1961 ynm ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1962 o zpm avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1963 a_30500_8700# zpp a_30200_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1964 a_23300_n3300# bna a_23000_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1965 a_27200_n3300# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1966 a_37400_100# znp a_37100_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1967 a_29000_6100# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1968 o znm a_72200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1969 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1970 a_25700_6100# zpp a_25400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1971 znm enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1972 ynp znp a_54800_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1973 a_64700_6100# zpp a_64400_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1974 a_22400_6100# zpp a_22100_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1975 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1976 a_59000_n1600# znp a_58700_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1977 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1978 a_29600_100# bna a_29300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1979 a_18200_7400# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1980 a_41000_10000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1981 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1982 avss bna a_21200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1983 a_57200_7400# bpa a_56900_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1984 avdd zpp a_44600_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1985 a_25400_n1600# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1986 a_48800_10000# zpp a_48500_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1987 a_29300_n1600# bna a_29000_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1988 a_47600_1800# bna a_47300_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1989 a_20000_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1990 avdd bpa a_20600_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1991 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1992 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1993 a_44300_1800# bnb a_44000_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1994 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1995 avdd bpa a_16400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1996 bpa_ bpa a_800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1997 a_55700_8700# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1998 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1999 a_9200_7400# bpa a_8900_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2000 a_52400_8700# bpa wp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2001 bpa_ bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2002 ynm znp a_66800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2003 bpb bpb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2004 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2005 a_7700_8700# bpa a_7400_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2006 ynp znp a_33200_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2007 a_44300_6100# zpp a_44000_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2008 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2009 a_37400_n3300# znp a_37100_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2010 a_16100_n3300# bna a_15800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2011 a_50900_100# znp a_50600_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2012 a_20000_n3300# bna a_19700_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2013 ypp zpp a_45800_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2014 a_69500_1800# znp a_69200_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2015 a_60200_100# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2016 a_27200_1800# ip ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2017 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2018 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2019 a_66200_1800# bnb zpm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2020 ynp im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2021 avss enb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2022 bna_ bnb a_6800_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2023 a_31700_n1600# znp a_31400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2024 zpm en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2025 a_55100_10000# bpb a_54800_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2026 a_35300_8700# bpa a_35000_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2027 a_35600_n1600# znp a_35300_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2028 wn bna a_42800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2029 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2030 avdd zpm o avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2031 a_39500_n1600# znp a_39200_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2032 avdd bpa a_21200_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2033 a_52400_100# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2034 a_25400_10000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2035 a_29300_10000# zpp a_29000_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2036 ypm zpp zpm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2037 a_27200_6100# zpp a_26900_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2038 zpm zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2039 a_44600_100# bnb a_44300_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2040 a_29000_7400# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2041 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2042 a_43700_n3300# bnb a_43400_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2043 a_11600_100# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2044 a_25700_7400# zpp a_25400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2045 a_47600_n3300# bna a_47300_n3300# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2046 a_64700_7400# zpp a_64400_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2047 a_16100_1800# bna a_15800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2048 a_22400_7400# zpp a_22100_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2049 a_69800_100# znp a_69500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2050 a_18200_8700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2051 ynp znp a_54800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2052 zpm bpb znm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2053 a_12800_1800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2054 a_57200_8700# bpa a_56900_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2055 a_36800_100# znp a_36500_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2056 a_51800_1800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2057 a_63200_n1600# bnb znm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2058 avdd bpa a_20600_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2059 a_41900_n1600# bna a_41600_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2060 bpa_ bpa a_800_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2061 a_45800_n1600# bnb a_45500_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2062 bna_ bnb a_6800_1800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2063 a_9200_8700# bpa a_8900_8700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2064 a_49700_n1600# znp a_49400_n1600# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2065 a_29000_100# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2066 a_3800_1800# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2067 a_16100_6100# bpa a_15800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2068 a_31700_10000# bpa a_31400_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2069 a_12200_n1600# bnb bna_ avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2070 a_55100_6100# bpb a_54800_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2071 a_35600_10000# bpa a_35300_10000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2072 bpa enb bpa_ avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2073 xp im ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2074 ynm znp a_38000_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2075 a_51800_6100# bpb a_51500_6100# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2076 zpp zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X2077 bnb bnb a_9800_100# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2078 a_3200_n1600# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2079 a_44300_7400# zpp a_44000_7400# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
.ends

.subckt sky130_rodovalho_ip__lpopamp im ip o ib en enb avdd vsub avss
Xslice0 im ip o en enb avdd avss bpa bpb bnb bna xp ypm ypp zpm zpp xn ynm ynp znm
+ znp vsub lpopamp_slice
Xslice1 im ip o en enb avdd avss bpa bpb bnb bna xp ypm ypp zpm zpp xn ynm ynp znm
+ znp vsub lpopamp_slice
X0 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X1 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X2 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X3 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X4 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X5 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X6 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X7 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X8 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X9 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X10 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X11 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X12 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X13 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X14 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X15 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X16 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X17 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X18 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X19 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X20 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=5.5
X21 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X22 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
X23 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
R0 ib bnb sky130_fd_pr__res_generic_m4 w=0.5 l=0.5
X24 ypm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=5.5
X25 ynm o sky130_fd_pr__cap_mim_m3_1 l=7.5 w=30
.ends

.subckt chipalooza_testchip1 gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12]
+ gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[1] gpio_analog[2]
+ gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6] gpio_analog[7] gpio_analog[8]
+ gpio_analog[9] gpio_noesd[0] gpio_noesd[10] gpio_noesd[11] gpio_noesd[12] gpio_noesd[13]
+ gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17] gpio_noesd[1] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6] gpio_noesd[7] gpio_noesd[8]
+ gpio_noesd[9] io_analog[0] io_analog[10] io_analog[1] io_analog[2] io_analog[3]
+ io_analog[4] io_analog[7] io_analog[8] io_analog[9] io_analog[5] io_analog[6] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24]
+ io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] vccd1 vccd2 vdda1 vdda2 m2_224722_800# m2_185716_800#
+ m2_35602_800# m3_800_35586# m2_128980_800# m2_522586_800# m2_572230_800# m2_106522_800#
+ m2_543862_800# m2_86428_800# m3_584320_272394# m2_58060_800# m3_800_508784# m2_29692_800#
+ m2_40330_800# m2_157348_800# m2_11962_800# m2_217630_800# sky130_ht_ip__hsxo_cpz1_0/power_gating_0/SG_AVSS
+ m2_111250_800# m2_178624_800# m2_28510_800# m3_800_466744# m3_584320_21256# m3_584320_7072#
+ m2_91156_800# m2_199900_800# m2_515494_800# m2_476488_800# m2_62788_800# m4_319794_703100#
+ m2_536770_800# m2_79336_800# m2_430390_800# m2_497764_800# m2_7234_800# m2_391384_800#
+ m2_61606_800# m4_176694_703100# m2_238906_800# m3_800_249652# m2_132526_800# m3_800_5890#
+ m2_565138_800# sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_1/vt m2_84064_800#
+ m2_153802_800# m2_469396_800# m2_480034_800# m2_55696_800# m3_584320_587908# m2_33238_800#
+ m2_451666_800# m2_76972_800# m2_384292_800# m2_4870_800# m2_54514_800# m3_584320_92372#
+ m2_472942_800# m3_327594_703100# m2_104158_800# m3_584320_452882# m2_125434_800#
+ m2_558046_800# m2_146710_800# m2_529678_800# m2_540316_800# m2_579322_800# m3_584320_12982#
+ m2_423298_800# m2_511948_800# m3_800_122030# m2_26146_800# m2_444574_800# m2_30874_800#
+ m2_69880_800# m3_800_335896# m2_47422_800# m2_465850_800# m2_101794_800# m4_228394_703100#
+ m2_584050_800# sky130_ajc_ip__por_0/por_ana_0/comparator_1/vt m2_118342_800# m3_800_293856#
+ m2_100612_800# m2_98248_800# m2_533224_800# m2_494218_800# m2_80518_800# m2_52150_800#
+ m2_504856_800# m2_554500_800# m2_19054_800# m2_437482_800# m2_23782_800# m3_584320_409642#
+ m2_398476_800# m3_800_14164# m2_123070_800# m2_292096_800# m2_380746_800# m2_22600_800#
+ m2_139618_800# m2_526132_800# m2_95884_800# m2_487126_800# m2_73426_800# m2_1324_800#
+ m5_319794_703100# m2_458758_800# m3_584320_497304# m2_16690_800# m2_94702_800# m4_166394_703100#
+ m2_352378_800# m2_412660_800# m2_581686_800# m2_373654_800# m2_115978_800# m5_176694_703100#
+ m2_394930_800# m3_171694_703100# m2_580504_800# m2_45058_800# m2_547408_800# m2_519040_800#
+ m2_88792_800# m2_441028_800# m2_66334_800# m2_501310_800# m2_462304_800# m2_37966_800#
+ m2_87610_800# m2_345286_800# m2_15508_800# m2_433936_800# sky130_ajc_ip__por_0/por_ana_0/comparator_0/vt
+ m2_366562_800# m2_108886_800# m3_800_423522# m3_584320_316816# m2_260182_800# m3_174194_703100#
+ m2_71062_800# m2_107704_800# m2_42694_800# m3_800_465562# m2_20236_800# m2_59242_800#
+ m2_63970_800# m2_405568_800# m3_584320_363220# m3_584320_454064# m3_800_4708# m2_455212_800#
+ m2_41512_800# sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_0/vt m3_800_79990#
+ m2_338194_800# m2_426844_800# m4_218094_703100# m2_299188_800# m2_320464_800# m2_387838_800#
+ m2_359470_800# m2_112432_800# m2_281458_800# m2_253090_800# m5_228394_703100# m2_341740_800#
+ m2_92338_800# sky130_be_ip__lsxo_0/dvss_ip m2_9598_800# m3_223394_703100# m3_800_337078#
+ m3_584320_3526# m2_13144_800# m2_8416_800# m2_448120_800# sky130_be_ip__lsxo_0/avss_ip
+ m2_34420_800# m2_370108_800# m3_584320_17710# m3_584320_586726# sky130_ht_ip__hsxo_cpz1_0/power_gating_0/EG_AVSS
+ m2_419752_800# m2_313372_800# m2_105340_800# m2_274366_800# m2_85246_800# m2_245998_800#
+ m2_295642_800# m2_56878_800# m3_584320_47714# m3_800_36768# m2_160894_800# m2_508402_800#
+ m2_10780_800# m4_330094_703100# m2_402022_800# m3_800_9436# m2_363016_800# m3_584320_362038#
+ m3_584320_273576# m5_166394_703100# m2_334648_800# m3_800_509966# m2_306280_800#
+ m2_267274_800# m2_355924_800# m2_78154_800# m2_82882_800# m2_288550_800# m2_6052_800#
+ m2_49786_800# m2_60424_800# m2_182170_800# m3_584320_22438# m2_99430_800# m3_800_292674#
+ m2_110068_800# m2_270820_800# m3_584320_8254# m2_27328_800# m2_81700_800# m2_48604_800#
+ m2_102976_800# m3_584320_16528# m2_327556_800# m3_584320_408460# m2_377200_800#
+ m2_119524_800# m2_221176_800# m2_348832_800# m2_32056_800# m2_242452_800# m2_75790_800#
+ m2_53332_800# m3_584320_498486# m2_24964_800# m2_416206_800# m2_124252_800# m2_561592_800#
+ m5_218094_703100# m2_331102_800# m3_800_10618# m3_584320_93554# m2_214084_800# m3_800_379118#
+ m2_3688_800# m2_302734_800# m2_175078_800# m3_325094_703100# m2_263728_800# m2_235360_800#
+ m2_74608_800# m2_196354_800# m2_46240_800# m2_206992_800# m2_2506_800# m2_167986_800#
+ m2_17872_800# m2_409114_800# m2_117160_800# m3_800_123212# m2_582868_800# m3_319794_703100#
+ m3_584320_317998# m2_97066_800# m2_324010_800# m2_68698_800# m3_584320_11800# m2_285004_800#
+ m3_176694_703100# m3_800_78808# m2_50968_800# m2_256636_800# m2_89974_800# m3_800_422340#
+ m2_150256_800# m2_67516_800# m2_189262_800# m2_277912_800# m2_121888_800# m2_171532_800#
+ m3_800_380300# m5_330094_703100# m2_575776_800# m2_120706_800# m3_800_15346# analog_mux_sel1v8_1/out
+ m2_228268_800# m2_72244_800# m2_490672_800# m2_316918_800# gpio_analog[17] m2_39148_800#
+ vssa2 m2_210538_800# m2_43876_800# m2_249544_800# m2_93520_800# m2_143164_800# m2_21418_800#
+ m2_231814_800# m3_225894_703100# m2_114796_800# m2_192808_800# m2_164440_800# m3_584320_2344#
+ m2_568684_800# m2_113614_800# m2_550954_800# m3_800_250834# vssd2 m2_65152_800#
+ m2_483580_800# m2_309826_800# m3_584320_48896# m2_203446_800# m2_36784_800# vssa1
+ m3_228394_703100# vssd1 m2_14326_800# m2_136072_800#
Xsky130_be_ip__lsxo_0 io_analog[3] vccd1 bias_generator_0/src_50 la_data_out[86] la_data_out[85]
+ io_out[12] gpio_noesd[4] gpio_noesd[3] sky130_be_ip__lsxo_0/avss_ip sky130_be_ip__lsxo_0/dvss_ip
+ vssa1 vssd1 sky130_be_ip__lsxo
Xbias_generator_0 gpio_analog[17] la_data_out[48] la_data_out[79] la_data_out[47]
+ bias_generator_0/src_10000_0 lpopamp_0/ib la_data_out[46] la_data_out[45] bias_generator_0/src_600
+ la_data_out[44] bias_generator_0/src_400 la_data_out[43] bias_generator_0/src_200_0
+ la_data_out[42] bias_generator_0/src_200_1 la_data_out[41] bias_generator_0/src_200_2
+ la_data_out[40] bias_generator_0/src_100 la_data_out[39] bias_generator_0/src_50
+ la_data_out[80] bias_generator_0/snk_2000 isolated_switch_ena1v8_2/in la_data_out[82]
+ bias_generator_0/snk_5000_2 bias_generator_0/snk_3700 la_data_out[83] la_data_out[78]
+ bias_generator_0/snk_test0 bias_generator_0/snk_test1 la_data_out[84] bias_generator_0/src_test1
+ la_data_out[38] analog_mux_sel1v8_5/inB la_data_out[49] bias_generator_0/snk_5000_0
+ la_data_out[125] vssd1 la_data_out[81] vdda1 vssa1 bias_generator
Xpower_stage_0[0] la_data_out[50] io_analog[5] vccd2 vccd2 vssd2 vssd2 power_stage
Xpower_stage_0[1] la_data_out[52] io_analog[6] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[2] la_data_out[54] io_analog[7] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[3] la_data_out[56] io_analog[8] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[4] la_data_out[58] io_analog[9] vccd2 vccd2 vssd2 vssd2 power_stage
Xpower_stage_0[5] la_data_out[60] io_analog[10] vdda2 vccd2 vssa2 vssd2 power_stage
Xpower_stage_0[6] la_data_out[62] power_stage_0[6]/sw_node vdda2 vccd2 vssa2 vssd2
+ power_stage
Xsky130_ajc_ip__overvoltage_0 io_analog[1] vccd1 analog_mux_sel1v8_0/inB io_out[6]
+ sky130_ajc_ip__overvoltage_0/itest la_data_out[105] la_data_out[104] la_data_out[103]
+ la_data_out[102] sky130_ajc_ip__overvoltage_0/vin la_data_out[100] la_data_out[101]
+ bias_generator_0/src_200_1 vssa1 vssd1 sky130_ajc_ip__overvoltage
Xsky130_ajc_ip__brownout_0 io_analog[0] io_out[0] vccd1 sky130_ajc_ip__brownout_0/osc_ck
+ io_out[1] analog_mux_sel1v8_0/inB la_data_out[112] la_data_out[113] la_data_out[111]
+ sky130_ajc_ip__brownout_0/itest sky130_ajc_ip__brownout_0/brout_filt la_data_out[107]
+ la_data_out[106] la_data_out[108] sky130_ajc_ip__brownout_0/vin_brout la_data_out[109]
+ la_data_out[115] sky130_ajc_ip__brownout_0/vin_vunder la_data_out[114] la_data_in[117]
+ io_out[5] la_data_out[116] la_data_out[110] bias_generator_0/src_200_0 sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_1/vt
+ sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_0/vt vssa1 vssd1 sky130_ajc_ip__brownout
Xpower_stage_1[0] la_data_out[77] io_analog[0] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[1] la_data_out[75] io_analog[1] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[2] la_data_out[73] io_analog[2] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[3] la_data_out[71] power_stage_1[3]/sw_node vdda1 vccd1 vssa1 vssd1
+ power_stage
Xpower_stage_1[4] la_data_out[69] io_analog[3] vdda1 vccd1 vssa1 vssd1 power_stage
Xpower_stage_1[5] la_data_out[67] power_stage_1[5]/sw_node vdda1 vccd1 vssa1 vssd1
+ power_stage
Xpower_stage_1[6] la_data_out[65] io_analog[4] vdda1 vccd1 vssa1 vssd1 power_stage
Xsky130_td_ip__opamp_hp_0 io_analog[10] gpio_noesd[7] bias_generator_0/src_100 analog_mux_sel1v8_1/inA
+ analog_mux_sel1v8_2/inA vccd2 la_data_out[37] vssd2 vssa2 sky130_td_ip__opamp_hp
Xanalog_mux_sel1v8_0 la_data_out[122] vccd1 gpio_noesd[2] analog_mux_sel1v8_0/inA
+ analog_mux_sel1v8_0/inB vdda1 vssa1 vssd1 analog_mux_sel1v8
Xanalog_mux_sel1v8_1 la_data_out[36] vccd2 analog_mux_sel1v8_1/out analog_mux_sel1v8_1/inA
+ analog_mux_sel1v8_1/inB vdda2 vssa2 vssd2 analog_mux_sel1v8
Xanalog_mux_sel1v8_2 la_data_out[34] vccd2 gpio_analog[9] analog_mux_sel1v8_2/inA
+ analog_mux_sel1v8_2/inB vdda2 vssa2 vssd2 analog_mux_sel1v8
Xanalog_mux_sel1v8_3 la_data_out[22] vccd2 gpio_analog[12] analog_mux_sel1v8_3/inA
+ lpopamp_0/ip vdda2 vssa2 vssd2 analog_mux_sel1v8
Xanalog_mux_sel1v8_4 la_data_out[23] vccd2 gpio_analog[11] analog_mux_sel1v8_4/inA
+ lpopamp_0/im vdda2 vssa2 vssd2 analog_mux_sel1v8
Xsky130_ht_ip__hsxo_cpz1_0 gpio_analog[15] gpio_analog[14] la_data_out[19] la_data_out[20]
+ io_out[23] io_analog[6] vccd2 vssd2 bias_generator_0/src_10000_0 sky130_ht_ip__hsxo_cpz1_0/power_gating_0/EG_AVSS
+ vssa2 vssd2 sky130_ht_ip__hsxo_cpz1_0/power_gating_0/SG_AVSS sky130_ht_ip__hsxo_cpz1
Xisolated_switch_ena1v8_0 la_data_out[123] vccd1 bias_generator_0/snk_3700 gpio_analog[5]
+ vdda1 vssd1 vssa1 isolated_switch_ena1v8
Xanalog_mux_sel1v8_5 la_data_out[18] vccd2 gpio_analog[16] analog_mux_sel1v8_5/inA
+ analog_mux_sel1v8_5/inB vdda2 vssa2 vssd2 analog_mux_sel1v8
Xisolated_switch_ena1v8_1 la_data_out[118] vccd1 bias_generator_0/snk_test0 gpio_analog[0]
+ vdda1 vssd1 vssa1 isolated_switch_ena1v8
Xisolated_switch_ena1v8_2 la_data_out[121] vccd1 isolated_switch_ena1v8_2/in gpio_analog[1]
+ vdda1 vssd1 vssa1 isolated_switch_ena1v8
Xsky130_vbl_ip__overvoltage_0 io_analog[4] vccd1 la_data_out[91] la_data_out[87] bias_generator_0/src_600
+ la_data_out[88] io_out[13] analog_mux_sel1v8_0/inA la_data_out[89] la_data_out[90]
+ vssd1 vssa1 sky130_vbl_ip__overvoltage
Xisolated_switch_ena1v8_4 la_data_out[124] vccd1 bias_generator_0/snk_test1 gpio_analog[6]
+ vdda1 vssd1 vssa1 isolated_switch_ena1v8
Xisolated_switch_ena1v8_5 la_data_out[17] vccd2 bias_generator_0/src_test1 gpio_analog[10]
+ vdda2 vssd2 vssa2 isolated_switch_ena1v8
Xlvl_shift_invert_0 la_data_out[21] vccd2 vdda2 lpopamp_0/enb lpopamp_0/en vssd2 lvl_shift_invert
Xsky130_od_ip__tempsensor_ext_vp_0 analog_mux_sel1v8_1/inB analog_mux_sel1v8_2/inB
+ la_data_out[35] analog_mux_sel1v8_0/inA io_analog[9] vssd2 sky130_od_ip__tempsensor_ext_vp
Xsky130_cw_ip__bandgap_0 la_data_out[1] la_data_out[3] la_data_out[4] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_data_out[10] la_data_out[11] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[2] analog_mux_sel1v8_5/inA
+ la_data_out[5] la_data_out[12] io_analog[5] vssd2 vssd2 sky130_cw_ip__bandgap
Xsky130_ajc_ip__por_0 io_analog[2] vccd1 analog_mux_sel1v8_0/inB la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[94] la_data_out[93] la_data_out[99] la_data_out[95]
+ bias_generator_0/src_200_2 sky130_ajc_ip__por_0/vin sky130_ajc_ip__por_0/porb_h
+ io_out[8] io_out[7] io_out[3] io_out[4] sky130_ajc_ip__por_0/itest la_data_in[120]
+ la_data_in[119] la_data_out[92] io_out[2] sky130_ajc_ip__por_0/por_ana_0/comparator_1/vt
+ sky130_ajc_ip__por_0/por_ana_0/comparator_0/vt vssa1 vssd1 sky130_ajc_ip__por
Xsky130_ak_ip__comparator_0 analog_mux_sel1v8_4/inA analog_mux_sel1v8_3/inA io_analog[8]
+ vssa2 la_data_out[28] la_data_out[29] la_data_out[30] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[33] la_data_out[32] la_data_out[31] io_out[17] vccd2
+ bias_generator_0/src_400 vssd2 sky130_ak_ip__comparator
Xlpopamp_0 lpopamp_0/im lpopamp_0/ip gpio_analog[13] lpopamp_0/ib lpopamp_0/en lpopamp_0/enb
+ io_analog[7] vssd2 vssa2 sky130_rodovalho_ip__lpopamp
R0 vssd1 io_oeb[13] sky130_fd_pr__res_generic_m3 w=0.56 l=0.7
R1 vssd1 io_oeb[5] sky130_fd_pr__res_generic_m3 w=0.335 l=0.435
R2 vssd1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.56 l=0.7
R3 io_oeb[17] vssd2 sky130_fd_pr__res_generic_m3 w=0.56 l=0.325
R4 vssd1 io_oeb[0] sky130_fd_pr__res_generic_m3 w=0.405 l=0.44
R5 vssd1 io_oeb[1] sky130_fd_pr__res_generic_m3 w=0.405 l=0.44
R6 io_oeb[23] vssd2 sky130_fd_pr__res_generic_m3 w=1.45 l=0.91
R7 vssd1 io_oeb[2] sky130_fd_pr__res_generic_m3 w=0.305 l=0.425
R8 vssd1 io_oeb[7] sky130_fd_pr__res_generic_m3 w=0.56 l=0.7
R9 vssd1 io_oeb[3] sky130_fd_pr__res_generic_m3 w=0.305 l=0.425
R10 vssd1 io_oeb[4] sky130_fd_pr__res_generic_m3 w=0.305 l=0.425
R11 vssd1 io_oeb[8] sky130_fd_pr__res_generic_m3 w=0.56 l=0.7
R12 vssd1 io_oeb[6] sky130_fd_pr__res_generic_m3 w=0.37 l=0.45
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xchipalooza_testchip1_0 gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12]
+ gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[1] gpio_analog[2]
+ gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6] gpio_analog[7] gpio_analog[8]
+ gpio_analog[9] gpio_noesd[0] gpio_noesd[10] gpio_noesd[11] gpio_noesd[12] gpio_noesd[13]
+ gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17] gpio_noesd[1] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6] gpio_noesd[7] gpio_noesd[8]
+ gpio_noesd[9] io_analog[0] io_analog[10] io_analog[1] io_analog[2] io_analog[3]
+ io_analog[4] io_analog[7] io_analog[8] io_analog[9] io_analog[5] io_analog[6] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24]
+ io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] vccd1 vccd2 vdda1 vdda2 la_oenb[27] la_oenb[16] wbs_dat_i[6]
+ io_in[23] la_oenb[0] la_oenb[111] la_oenb[125] wbs_dat_i[26] la_oenb[117] wbs_dat_o[20]
+ io_in_3v3[7] wbs_dat_o[12] io_in[14] wbs_dat_o[4] wbs_dat_o[7] la_oenb[8] wbs_sel_i[0]
+ la_oenb[25] chipalooza_testchip1_0/sky130_ht_ip__hsxo_cpz1_0/power_gating_0/SG_AVSS
+ wbs_dat_o[27] la_oenb[14] wbs_dat_i[4] io_in_3v3[15] io_in_3v3[4] io_in_3v3[1] wbs_adr_i[22]
+ la_oenb[20] la_oenb[109] la_oenb[98] wbs_adr_i[14] io_analog[4] la_oenb[115] wbs_dat_o[18]
+ la_oenb[85] la_oenb[104] wbs_we_i la_oenb[74] wbs_dat_o[13] io_analog[6] la_oenb[31]
+ io_in[20] la_oenb[1] io_in_3v3[26] la_oenb[123] chipalooza_testchip1_0/sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_1/vt
+ wbs_adr_i[20] la_oenb[7] la_oenb[96] la_oenb[99] wbs_adr_i[12] io_in[13] wbs_dat_o[5]
+ la_oenb[91] wbs_adr_i[18] la_oenb[72] wbs_cyc_i wbs_dat_o[11] io_in_3v3[6] la_oenb[97]
+ io_clamp_high[0] wbs_dat_o[25] io_in_3v3[11] wbs_dat_o[31] la_oenb[121] la_oenb[5]
+ la_oenb[113] la_oenb[116] la_oenb[127] io_in[2] la_oenb[83] la_oenb[108] io_in[21]
+ wbs_sel_i[3] la_oenb[89] wbs_adr_i[5] wbs_adr_i[16] io_in[18] wbs_dat_o[9] la_oenb[95]
+ wbs_adr_i[25] io_analog[5] user_irq[2] chipalooza_testchip1_0/sky130_ajc_ip__por_0/por_ana_0/comparator_1/vt
+ wbs_dat_o[29] io_in_3v3[19] wbs_dat_o[24] wbs_adr_i[24] la_oenb[114] la_oenb[103]
+ wbs_adr_i[19] wbs_adr_i[11] la_oenb[106] la_oenb[120] wbs_dat_i[2] la_oenb[87] wbs_dat_i[3]
+ io_in[10] la_oenb[76] io_in[24] wbs_adr_i[31] la_oenb[46] la_oenb[71] wbs_adr_i[3]
+ la_oenb[3] la_oenb[112] wbs_dat_i[23] la_oenb[101] wbs_adr_i[17] wb_clk_i io_analog[4]
+ la_oenb[93] io_in_3v3[12] wbs_sel_i[1] wbs_adr_i[23] io_analog[6] la_oenb[63] la_oenb[80]
+ user_irq[0] la_oenb[69] wbs_adr_i[29] io_analog[6] la_oenb[75] io_clamp_low[2] user_clock2
+ wbs_adr_i[9] la_oenb[118] la_oenb[110] wbs_dat_i[21] la_oenb[88] wbs_adr_i[15] la_oenb[105]
+ la_oenb[94] wbs_adr_i[7] wbs_adr_i[21] la_oenb[61] wbs_dat_o[1] la_oenb[86] chipalooza_testchip1_0/sky130_ajc_ip__por_0/por_ana_0/comparator_0/vt
+ la_oenb[67] wbs_adr_i[27] io_in_3v3[16] io_in_3v3[8] la_oenb[37] io_clamp_high[2]
+ wbs_dat_i[16] wbs_dat_o[26] wbs_dat_i[8] io_in[15] wbs_dat_o[2] wbs_adr_i[13] wbs_dat_i[14]
+ la_oenb[78] io_in[9] io_in[11] io_in[26] la_oenb[92] wbs_adr_i[8] chipalooza_testchip1_0/sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_0/vt
+ io_in_3v3[22] la_oenb[59] la_oenb[84] io_analog[5] la_oenb[48] la_oenb[54] la_oenb[73]
+ la_oenb[65] wbs_adr_i[28] la_oenb[43] la_oenb[35] io_analog[5] la_oenb[60] wbs_dat_i[22]
+ chipalooza_testchip1_0/sky130_be_ip__lsxo_0/dvss_ip wbs_dat_i[0] io_clamp_low[1]
+ io_in_3v3[18] io_in[0] wbs_adr_i[1] wbs_adr_i[0] la_oenb[90] chipalooza_testchip1_0/sky130_be_ip__lsxo_0/avss_ip
+ wbs_adr_i[6] la_oenb[68] io_in[3] io_in_3v3[13] chipalooza_testchip1_0/sky130_ht_ip__hsxo_cpz1_0/power_gating_0/EG_AVSS
+ la_oenb[82] la_oenb[52] wbs_adr_i[26] la_oenb[41] wbs_dat_i[20] la_oenb[33] la_oenb[47]
+ wbs_dat_i[12] io_in_3v3[5] io_in_3v3[23] la_oenb[9] la_oenb[107] wbs_dat_o[0] io_analog[4]
+ la_oenb[77] io_in[25] la_oenb[66] io_in_3v3[9] io_in[7] io_analog[6] la_oenb[58]
+ io_in_3v3[14] la_oenb[50] la_oenb[39] la_oenb[64] wbs_dat_i[18] wbs_dat_o[19] la_oenb[45]
+ wbs_stb_i wbs_dat_i[10] wbs_dat_i[13] la_oenb[15] io_in[4] wbs_dat_i[24] io_in[19]
+ wbs_dat_i[27] la_oenb[40] io_in[1] wbs_adr_i[4] wbs_dat_i[19] wbs_adr_i[10] wbs_dat_i[25]
+ io_in_3v3[3] la_oenb[56] io_in_3v3[10] la_oenb[70] wbs_adr_i[30] la_oenb[26] la_oenb[62]
+ wbs_dat_i[5] la_oenb[32] wbs_dat_o[17] wbs_dat_i[11] io_in[12] wbs_dat_o[3] la_oenb[81]
+ wbs_dat_i[31] la_oenb[122] io_analog[5] la_oenb[57] io_in_3v3[25] io_in[6] la_oenb[24]
+ io_in[17] wbs_ack_o la_oenb[49] la_oenb[13] io_clamp_low[0] la_oenb[38] la_oenb[30]
+ wbs_dat_i[17] la_oenb[19] wbs_dat_i[9] la_oenb[22] wb_rst_i la_oenb[11] wbs_adr_i[2]
+ la_oenb[79] wbs_dat_i[29] io_in_3v3[21] user_irq[1] io_analog[4] io_in[8] wbs_dat_o[23]
+ la_oenb[55] wbs_dat_o[15] io_in_3v3[2] la_oenb[44] io_analog[6] io_in[22] wbs_dat_o[10]
+ la_oenb[36] wbs_dat_o[21] io_in[16] la_oenb[6] wbs_dat_i[15] la_oenb[17] la_oenb[42]
+ wbs_dat_o[30] la_oenb[12] io_in_3v3[17] io_analog[4] la_oenb[126] wbs_dat_i[30]
+ io_in_3v3[24] gpio_analog[8] la_oenb[28] wbs_dat_o[16] la_oenb[102] la_oenb[53]
+ gpio_analog[17] wbs_dat_i[7] vssa2 la_oenb[23] wbs_dat_o[8] la_oenb[34] wbs_dat_o[22]
+ la_oenb[4] wbs_sel_i[2] la_oenb[29] io_clamp_high[1] wbs_dat_o[28] la_oenb[18] la_oenb[10]
+ io_in_3v3[0] la_oenb[124] wbs_dat_i[28] la_oenb[119] io_in_3v3[20] vssd2 wbs_dat_o[14]
+ la_oenb[100] la_oenb[51] io_in[5] la_oenb[21] wbs_dat_o[6] vssa1 io_analog[5] vssd1
+ wbs_dat_i[1] la_oenb[2] chipalooza_testchip1
.ends

