magic
tech sky130A
magscale 1 2
timestamp 1713926953
<< locali >>
rect 1990 -3266 2210 -2972
rect 2470 -3022 2519 -2972
rect 2470 -3215 2480 -3022
rect 2514 -3215 2519 -3022
rect 2470 -3266 2519 -3215
<< viali >>
rect 2480 -3215 2514 -3022
<< metal1 >>
rect 2062 294 2641 302
rect 2062 234 2122 294
rect 2063 216 2122 234
rect 2588 216 2641 294
rect 2063 154 2641 216
rect 2063 -2676 2115 154
rect 2150 -1558 2214 8
rect 2326 -654 2378 92
rect 2482 14 2641 154
rect 2470 -582 2641 14
rect 2326 -656 2374 -654
rect 2326 -674 2378 -662
rect 2326 -868 2378 -860
rect 2324 -922 2372 -920
rect 2324 -1666 2376 -922
rect 2324 -1668 2378 -1666
rect 2326 -1676 2378 -1668
rect 2326 -1870 2378 -1862
rect 2330 -1920 2380 -1918
rect 2063 -2818 2115 -2812
rect 2144 -3709 2208 -1990
rect 2144 -3967 2208 -3941
rect 2330 -3402 2384 -1920
rect 2480 -2574 2544 -1008
rect 2589 -2676 2641 -582
rect 2589 -2821 2641 -2812
rect 2470 -3001 2540 -2972
rect 2470 -3265 2540 -3239
rect 2330 -3967 2384 -3634
<< via1 >>
rect 2122 216 2588 294
rect 2326 -860 2378 -674
rect 2326 -1862 2378 -1676
rect 2063 -2812 2115 -2676
rect 2144 -3941 2208 -3709
rect 2589 -2812 2641 -2676
rect 2470 -3022 2540 -3001
rect 2470 -3215 2480 -3022
rect 2480 -3215 2514 -3022
rect 2514 -3215 2540 -3022
rect 2470 -3239 2540 -3215
rect 2330 -3634 2384 -3402
<< metal2 >>
rect 1990 294 2710 388
rect 1990 216 2122 294
rect 2588 216 2710 294
rect 1990 154 2710 216
rect 1990 -674 2710 -666
rect 1990 -860 2326 -674
rect 2378 -860 2710 -674
rect 1990 -900 2710 -860
rect 1990 -1676 2710 -1670
rect 1990 -1862 2326 -1676
rect 2378 -1862 2710 -1676
rect 1990 -1904 2710 -1862
rect 1990 -2676 2710 -2670
rect 1990 -2812 2063 -2676
rect 2115 -2812 2589 -2676
rect 2641 -2812 2710 -2676
rect 1990 -2904 2710 -2812
rect 1990 -3239 2470 -3001
rect 2540 -3239 2710 -3001
rect 2324 -3634 2330 -3402
rect 2384 -3634 2390 -3402
rect 2138 -3941 2144 -3709
rect 2208 -3941 2214 -3709
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ#1  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 ../../chipalooza/sky130_od_ip__tempsensor/mag
timestamp 1713474431
transform 1 0 2357 0 1 -3119
box -183 -183 183 183
use sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ  sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ_0
timestamp 1713888873
transform 1 0 2352 0 1 -2289
box -358 -597 358 597
use sky130_fd_pr__pfet_g5v0d10v5_H75TTW  sky130_fd_pr__pfet_g5v0d10v5_H75TTW_0
timestamp 1713888873
transform 1 0 2352 0 1 -281
box -358 -597 358 597
use sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ  XM13
timestamp 1713888873
transform 1 0 2352 0 1 -1285
box -358 -597 358 597
<< end >>
