magic
tech sky130A
magscale 1 2
timestamp 1713983242
<< psubdiff >>
rect 3348 5238 3808 5296
rect 3348 3328 3402 5238
rect 3750 3328 3808 5238
rect 3348 3288 3808 3328
<< psubdiffcont >>
rect 3402 3328 3750 5238
<< locali >>
rect 2942 6450 3028 6470
rect 2942 6126 2952 6450
rect 3016 6126 3028 6450
rect 2942 6112 3028 6126
rect 1184 5502 1430 5506
rect 1184 5374 1202 5502
rect 1410 5374 1430 5502
rect 1184 5366 1430 5374
rect 3340 5238 3794 5286
rect 3340 5074 3402 5238
rect 886 4922 3402 5074
rect 160 4712 3046 4722
rect 160 4638 166 4712
rect 3036 4638 3046 4712
rect 160 4632 3046 4638
rect 3340 3328 3402 4922
rect 3750 3328 3794 5238
rect 3340 3294 3794 3328
<< viali >>
rect 2952 6126 3016 6450
rect 1202 5374 1410 5502
rect 166 4638 3036 4712
<< metal1 >>
rect 896 6718 3020 6722
rect 558 6590 3020 6718
rect 558 6566 1128 6590
rect 558 5182 816 6566
rect 2942 6460 3174 6470
rect 2942 6450 3090 6460
rect 2942 6126 2952 6450
rect 3016 6126 3090 6450
rect 2942 6122 3090 6126
rect 3158 6122 3174 6460
rect 2942 6112 3174 6122
rect 896 5760 3500 6004
rect 908 5694 2994 5710
rect 908 5642 948 5694
rect 2938 5642 2994 5694
rect 908 5630 2994 5642
rect 1184 5502 1430 5508
rect 1184 5374 1202 5502
rect 1410 5374 1430 5502
rect 1184 5366 1430 5374
rect 558 5176 1004 5182
rect 16 4890 3012 5176
rect 3218 4742 3500 5760
rect 76 4712 3500 4742
rect 76 4638 166 4712
rect 3036 4638 3500 4712
rect 76 4530 3500 4638
rect 24 2544 234 2820
rect 3218 2780 3500 4530
rect 3944 2132 4146 2338
rect 12 1542 216 1750
rect 26 206 260 442
<< via1 >>
rect 3090 6122 3158 6460
rect 948 5642 2938 5694
rect 1202 5374 1410 5502
<< metal2 >>
rect 3082 6460 3168 6470
rect 3082 6122 3090 6460
rect 3158 6122 3168 6460
rect 40 5918 350 5924
rect 40 5694 2994 5918
rect 40 5642 948 5694
rect 2938 5642 2994 5694
rect 40 5614 2994 5642
rect 1184 5502 1430 5508
rect 30 5494 230 5498
rect 1184 5494 1202 5502
rect 30 5374 1202 5494
rect 1410 5374 1430 5502
rect 30 5372 1430 5374
rect 30 5298 230 5372
rect 1184 5366 1430 5372
rect 3082 3530 3168 6122
rect 1632 3478 3168 3530
use isolated_switch  isolated_switch_0
timestamp 1713983242
transform 1 0 -301 0 1 2911
box 301 -2911 4463 1830
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 896 0 1 5065
box -66 -43 2178 1671
<< labels >>
flabel metal1 16 4890 348 5176 0 FreeSans 560 0 0 0 dvss
port 0 nsew
flabel metal2 30 5298 230 5498 0 FreeSans 560 0 0 0 on
port 1 nsew
flabel metal2 40 5614 350 5924 0 FreeSans 560 0 0 0 dvdd
port 2 nsew
flabel metal1 12 1542 216 1750 0 FreeSans 560 0 0 0 in
port 3 nsew
flabel metal1 24 2544 234 2820 0 FreeSans 560 0 0 0 avdd
port 4 nsew
flabel metal1 26 206 260 442 0 FreeSans 560 0 0 0 avss
port 5 nsew
flabel metal1 3944 2132 4146 2338 0 FreeSans 560 0 0 0 out
port 6 nsew
<< end >>
