* NGSPICE file created from bias_generator.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ a_n158_n300# a_n100_n388# a_100_n300#
+ a_n292_n522#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n292_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RK a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_QRKT8P a_n158_n300# a_n100_n388# a_100_n300# a_n292_n522#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n292_n522# sky130_fd_pr__nfet_05v0_nvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P a_n158_n300# a_n100_n388# a_100_n300#
+ a_n292_n522#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n292_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_nstack itail ena nbias avss vcasc
XXM12 avss nbias m1_3726_n2502# avss sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RK
XXM6 vcasc nbias m1_3726_n2502# avss sky130_fd_pr__nfet_05v0_nvt_QRKT8P
XXM7 vcasc ena itail avss sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P
.ends

.subckt sky130_fd_pr__res_high_po_0p35_P35QVK a_380_2984# a_5692_n3416# a_n3770_2984#
+ a_3866_2984# a_3202_n3416# a_n1446_n3416# a_n284_n3416# a_n616_2984# a_4696_n3416#
+ a_4198_2984# a_2206_n3416# a_n1114_2984# a_n4102_2984# a_n616_n3416# a_6190_n3416#
+ a_n6592_2984# a_2372_2984# a_n5762_n3416# a_5360_2984# a_214_2984# a_n3604_2984#
+ a_1210_n3416# a_5194_n3416# a_6522_n3416# a_n4766_n3416# a_1874_2984# a_4862_2984#
+ a_4198_n3416# a_5526_n3416# a_5194_2984# a_n6260_n3416# a_878_n3416# a_n3438_2984#
+ a_n2110_2984# a_n6426_2984# a_2206_2984# a_n118_n3416# a_n3770_n3416# a_4696_2984#
+ a_n5264_n3416# a_48_2984# a_4530_n3416# a_n2774_n3416# a_n1612_2984# a_n4600_2984#
+ a_n5928_2984# a_1708_2984# a_6024_n3416# a_n4268_n3416# a_2870_2984# a_3534_n3416#
+ a_712_2984# a_n1778_n3416# a_5028_2984# a_5028_n3416# a_n948_2984# a_2538_n3416#
+ a_6190_2984# a_n1446_2984# a_n3272_n3416# a_n4434_2984# a_n4600_n3416# a_3202_2984#
+ a_n948_n3416# a_5692_2984# a_380_n3416# a_546_2984# a_4032_n3416# a_n2276_n3416#
+ a_n3604_n3416# a_n3936_2984# a_1542_n3416# a_2704_2984# a_3036_n3416# a_712_n3416#
+ a_n2608_n3416# a_n4268_2984# a_3036_2984# a_6024_2984# a_5858_n3416# a_n1280_n3416#
+ a_n6592_n3416# a_n2442_2984# a_n4102_n3416# a_2538_2984# a_n5430_2984# a_2040_n3416#
+ a_5526_2984# a_1210_2984# a_n1612_n3416# a_n5596_n3416# a_4862_n3416# a_n450_n3416#
+ a_n1944_2984# a_n3106_n3416# a_n4932_2984# a_1044_n3416# a_n450_2984# a_3700_2984#
+ a_6356_n3416# a_214_n3416# a_n5928_n3416# a_n6722_n3546# a_3866_n3416# a_n2276_2984#
+ a_n5264_2984# a_1044_2984# a_4032_2984# a_n2110_n3416# a_n6094_n3416# a_n1778_2984#
+ a_n4766_2984# a_5360_n3416# a_n284_2984# a_3534_2984# a_n4932_n3416# a_6522_2984#
+ a_n1114_n3416# a_2870_n3416# a_n5098_n3416# a_n6426_n3416# a_878_2984# a_4364_n3416#
+ a_n5098_2984# a_n3936_n3416# a_n2940_2984# a_1874_n3416# a_3368_n3416# a_n3272_2984#
+ a_3368_2984# a_48_n3416# a_n6260_2984# a_2040_2984# a_6356_2984# a_n5430_n3416#
+ a_n2940_n3416# a_n118_2984# a_n2774_2984# a_n4434_n3416# a_n5762_2984# a_1542_2984#
+ a_2372_n3416# a_4530_2984# a_5858_2984# a_3700_n3416# a_n1944_n3416# a_n3438_n3416#
+ a_n6094_2984# a_n782_n3416# a_1376_n3416# a_n782_2984# a_2704_n3416# a_546_n3416#
+ a_n3106_2984# a_n1280_2984# a_n5596_2984# a_1376_2984# a_1708_n3416# a_4364_2984#
+ a_n2442_n3416# a_n2608_2984#
X0 a_n3936_2984# a_n3936_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X1 a_n1612_2984# a_n1612_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X2 a_n6592_2984# a_n6592_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X3 a_n4434_2984# a_n4434_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X4 a_48_2984# a_48_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X5 a_2704_2984# a_2704_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X6 a_4862_2984# a_4862_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X7 a_3202_2984# a_3202_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X8 a_5360_2984# a_5360_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X9 a_5526_2984# a_5526_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X10 a_n948_2984# a_n948_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X11 a_n782_2984# a_n782_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X12 a_6024_2984# a_6024_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X13 a_n4932_2984# a_n4932_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X14 a_1376_2984# a_1376_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X15 a_878_2984# a_878_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X16 a_4198_2984# a_4198_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X17 a_n3770_2984# a_n3770_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X18 a_n1446_2984# a_n1446_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X19 a_3700_2984# a_3700_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X20 a_n4268_2984# a_n4268_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X21 a_n2110_2984# a_n2110_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X22 a_1874_2984# a_1874_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X23 a_6522_2984# a_6522_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X24 a_2372_2984# a_2372_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X25 a_2538_2984# a_2538_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X26 a_4696_2984# a_4696_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X27 a_3036_2984# a_3036_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X28 a_5194_2984# a_5194_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X29 a_n1944_2984# a_n1944_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X30 a_n4766_2984# a_n4766_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X31 a_n2608_2984# a_n2608_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X32 a_n2442_2984# a_n2442_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X33 a_214_2984# a_214_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X34 a_n5430_2984# a_n5430_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X35 a_n5264_2984# a_n5264_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X36 a_n3106_2984# a_n3106_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X37 a_2870_2984# a_2870_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X38 a_n1280_2984# a_n1280_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X39 a_1210_2984# a_1210_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X40 a_3534_2984# a_3534_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X41 a_5692_2984# a_5692_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X42 a_5858_2984# a_5858_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X43 a_712_2984# a_712_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X44 a_4032_2984# a_4032_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X45 a_6190_2984# a_6190_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X46 a_6356_2984# a_6356_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X47 a_n5928_2984# a_n5928_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X48 a_n5762_2984# a_n5762_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X49 a_n3604_2984# a_n3604_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X50 a_n118_2984# a_n118_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X51 a_n6426_2984# a_n6426_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X52 a_n4102_2984# a_n4102_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X53 a_n1778_2984# a_n1778_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X54 a_4530_2984# a_4530_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X55 a_n4600_2984# a_n4600_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X56 a_n2276_2984# a_n2276_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X57 a_n5098_2984# a_n5098_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X58 a_n616_2984# a_n616_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X59 a_1044_2984# a_1044_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X60 a_3368_2984# a_3368_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X61 a_546_2984# a_546_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X62 a_n2940_2984# a_n2940_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X63 a_n2774_2984# a_n2774_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X64 a_380_2984# a_380_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X65 a_n5596_2984# a_n5596_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X66 a_n3438_2984# a_n3438_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X67 a_n3272_2984# a_n3272_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X68 a_n1114_2984# a_n1114_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X69 a_n6260_2984# a_n6260_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X70 a_n6094_2984# a_n6094_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X71 a_1708_2984# a_1708_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X72 a_1542_2984# a_1542_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X73 a_2206_2984# a_2206_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X74 a_3866_2984# a_3866_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X75 a_2040_2984# a_2040_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X76 a_4364_2984# a_4364_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X77 a_5028_2984# a_5028_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X78 a_n450_2984# a_n450_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X79 a_n284_2984# a_n284_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ w_n358_n597# a_n158_n300# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n358_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_H75TTW w_n358_n597# a_n158_n300# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n358_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_pstack avdd avss pcasc enb itail vcasc pbias
XXM13 avdd m1_2150_n1558# pcasc vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__pfet_g5v0d10v5_G8LMTZ_0 avdd itail enb vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss enb sky130_fd_pr__diode_pw2nd_05v5_FT76RK
Xsky130_fd_pr__pfet_g5v0d10v5_H75TTW_0 avdd m1_2150_n1558# pbias avdd sky130_fd_pr__pfet_g5v0d10v5_H75TTW
.ends

.subckt bias_generator ref_in enb ena avss enb_10000_0 src_10000_0 src_10000_1 enb_10000_1
+ enb_600 src_600 enb_400 src_400 enb_200_0 src_200_0 enb_200_1 src_200_1 enb_200_2
+ src_200_2 enb_100 src_100 enb_50 src_50 ena_5000_0 snk_2000 ena_5000_1 snk_5000_1
+ ena_5000_2 snk_5000_2 snk_3700 ena_3700 ena_test0 snk_test0 snk_test1 ena_test1
+ src_test1 enb_test1 src_test0 enb_test0 avdd snk_5000_0 ena_2000
Xbias_nstack_0[0] snk_test0 ena_test0 bias_nstack_0[9]/nbias avss bias_nstack_0[0]/vcasc
+ bias_nstack
Xbias_nstack_0[1] snk_test0 ena_test0 bias_nstack_0[9]/nbias avss bias_nstack_0[1]/vcasc
+ bias_nstack
Xbias_nstack_0[2] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[2]/vcasc
+ bias_nstack
Xbias_nstack_0[3] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[3]/vcasc
+ bias_nstack
Xbias_nstack_0[4] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[4]/vcasc
+ bias_nstack
Xbias_nstack_0[5] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[5]/vcasc
+ bias_nstack
Xbias_nstack_0[6] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[6]/vcasc
+ bias_nstack
Xbias_nstack_0[7] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[7]/vcasc
+ bias_nstack
Xbias_nstack_0[8] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[8]/vcasc
+ bias_nstack
Xbias_nstack_0[9] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[9]/vcasc
+ bias_nstack
Xbias_nstack_0[10] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[10]/vcasc
+ bias_nstack
Xbias_nstack_0[11] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[11]/vcasc
+ bias_nstack
Xbias_nstack_0[12] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[12]/vcasc
+ bias_nstack
Xbias_nstack_0[13] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[13]/vcasc
+ bias_nstack
Xbias_nstack_0[14] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[14]/vcasc
+ bias_nstack
Xbias_nstack_0[15] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[15]/vcasc
+ bias_nstack
Xbias_nstack_0[16] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[16]/vcasc
+ bias_nstack
Xbias_nstack_0[17] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[17]/vcasc
+ bias_nstack
Xbias_nstack_0[18] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[18]/vcasc
+ bias_nstack
Xbias_nstack_0[19] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[19]/vcasc
+ bias_nstack
Xbias_nstack_0[20] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[20]/vcasc
+ bias_nstack
Xbias_nstack_0[21] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[21]/vcasc
+ bias_nstack
Xbias_nstack_0[22] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[22]/vcasc
+ bias_nstack
Xbias_nstack_0[23] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[23]/vcasc
+ bias_nstack
Xbias_nstack_0[24] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[24]/vcasc
+ bias_nstack
Xbias_nstack_0[25] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[25]/vcasc
+ bias_nstack
Xbias_nstack_0[26] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[26]/vcasc
+ bias_nstack
Xbias_nstack_0[27] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[27]/vcasc
+ bias_nstack
Xbias_nstack_0[28] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[28]/vcasc
+ bias_nstack
Xbias_nstack_0[29] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[29]/vcasc
+ bias_nstack
Xbias_nstack_0[30] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[30]/vcasc
+ bias_nstack
Xbias_nstack_0[31] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[31]/vcasc
+ bias_nstack
Xbias_nstack_0[32] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[32]/vcasc
+ bias_nstack
Xbias_nstack_0[33] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[33]/vcasc
+ bias_nstack
Xbias_nstack_0[34] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[34]/vcasc
+ bias_nstack
Xbias_nstack_0[35] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[35]/vcasc
+ bias_nstack
Xbias_nstack_0[36] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[36]/vcasc
+ bias_nstack
Xbias_nstack_0[37] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[37]/vcasc
+ bias_nstack
Xbias_nstack_0[38] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[38]/vcasc
+ bias_nstack
Xbias_nstack_0[39] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[39]/vcasc
+ bias_nstack
Xbias_nstack_0[40] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[40]/vcasc
+ bias_nstack
Xbias_nstack_0[41] snk_2000 ena_2000 bias_nstack_0[9]/nbias avss bias_nstack_0[41]/vcasc
+ bias_nstack
Xbias_nstack_0[42] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[43] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[44] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[45] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[46] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[47] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[48] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[49] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[50] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[51] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[52] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[53] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[54] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[55] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[56] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[57] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[58] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[59] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[60] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[61] bias_nstack_0[61]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[9]/nbias
+ bias_nstack
Xbias_nstack_0[62] bias_pstack_0[62]/itail ena bias_nstack_0[9]/nbias avss bias_nstack_0[62]/vcasc
+ bias_nstack
Xbias_nstack_0[63] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[63]/vcasc
+ bias_nstack
Xbias_nstack_0[64] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[64]/vcasc
+ bias_nstack
Xbias_nstack_0[65] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[65]/vcasc
+ bias_nstack
Xbias_nstack_0[66] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[66]/vcasc
+ bias_nstack
Xbias_nstack_0[67] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[67]/vcasc
+ bias_nstack
Xbias_nstack_0[68] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[68]/vcasc
+ bias_nstack
Xbias_nstack_0[69] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[69]/vcasc
+ bias_nstack
Xbias_nstack_0[70] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[70]/vcasc
+ bias_nstack
Xbias_nstack_0[71] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[71]/vcasc
+ bias_nstack
Xbias_nstack_0[72] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[72]/vcasc
+ bias_nstack
Xbias_nstack_0[73] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[73]/vcasc
+ bias_nstack
Xbias_nstack_0[74] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[74]/vcasc
+ bias_nstack
Xbias_nstack_0[75] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[75]/vcasc
+ bias_nstack
Xbias_nstack_0[76] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[76]/vcasc
+ bias_nstack
Xbias_nstack_0[77] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[77]/vcasc
+ bias_nstack
Xbias_nstack_0[78] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[78]/vcasc
+ bias_nstack
Xbias_nstack_0[79] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[79]/vcasc
+ bias_nstack
Xbias_nstack_0[80] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[80]/vcasc
+ bias_nstack
Xbias_nstack_0[81] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[81]/vcasc
+ bias_nstack
Xbias_nstack_0[82] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[82]/vcasc
+ bias_nstack
Xbias_nstack_0[83] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[83]/vcasc
+ bias_nstack
Xbias_nstack_0[84] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[84]/vcasc
+ bias_nstack
Xbias_nstack_0[85] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[85]/vcasc
+ bias_nstack
Xbias_nstack_0[86] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[86]/vcasc
+ bias_nstack
Xbias_nstack_0[87] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[87]/vcasc
+ bias_nstack
Xbias_nstack_0[88] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[88]/vcasc
+ bias_nstack
Xbias_nstack_0[89] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[89]/vcasc
+ bias_nstack
Xbias_nstack_0[90] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[90]/vcasc
+ bias_nstack
Xbias_nstack_0[91] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[91]/vcasc
+ bias_nstack
Xbias_nstack_0[92] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[92]/vcasc
+ bias_nstack
Xbias_nstack_0[93] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[93]/vcasc
+ bias_nstack
Xbias_nstack_0[94] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[94]/vcasc
+ bias_nstack
Xbias_nstack_0[95] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[95]/vcasc
+ bias_nstack
Xbias_nstack_0[96] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[96]/vcasc
+ bias_nstack
Xbias_nstack_0[97] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[97]/vcasc
+ bias_nstack
Xbias_nstack_0[98] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[98]/vcasc
+ bias_nstack
Xbias_nstack_0[99] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[99]/vcasc
+ bias_nstack
Xbias_nstack_0[100] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[100]/vcasc
+ bias_nstack
Xbias_nstack_0[101] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[101]/vcasc
+ bias_nstack
Xbias_nstack_0[102] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[102]/vcasc
+ bias_nstack
Xbias_nstack_0[103] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[103]/vcasc
+ bias_nstack
Xbias_nstack_0[104] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[104]/vcasc
+ bias_nstack
Xbias_nstack_0[105] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[105]/vcasc
+ bias_nstack
Xbias_nstack_0[106] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[106]/vcasc
+ bias_nstack
Xbias_nstack_0[107] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[107]/vcasc
+ bias_nstack
Xbias_nstack_0[108] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[108]/vcasc
+ bias_nstack
Xbias_nstack_0[109] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[109]/vcasc
+ bias_nstack
Xbias_nstack_0[110] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[110]/vcasc
+ bias_nstack
Xbias_nstack_0[111] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[111]/vcasc
+ bias_nstack
Xbias_nstack_0[112] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[112]/vcasc
+ bias_nstack
Xbias_nstack_0[113] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[113]/vcasc
+ bias_nstack
Xbias_nstack_0[114] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[114]/vcasc
+ bias_nstack
Xbias_nstack_0[115] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[115]/vcasc
+ bias_nstack
Xbias_nstack_0[116] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[116]/vcasc
+ bias_nstack
Xbias_nstack_0[117] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[117]/vcasc
+ bias_nstack
Xbias_nstack_0[118] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[118]/vcasc
+ bias_nstack
Xbias_nstack_0[119] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[119]/vcasc
+ bias_nstack
Xbias_nstack_0[120] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[120]/vcasc
+ bias_nstack
Xbias_nstack_0[121] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[121]/vcasc
+ bias_nstack
Xbias_nstack_0[122] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[122]/vcasc
+ bias_nstack
Xbias_nstack_0[123] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[123]/vcasc
+ bias_nstack
Xbias_nstack_0[124] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[124]/vcasc
+ bias_nstack
Xbias_nstack_0[125] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[125]/vcasc
+ bias_nstack
Xbias_nstack_0[126] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[126]/vcasc
+ bias_nstack
Xbias_nstack_0[127] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[127]/vcasc
+ bias_nstack
Xbias_nstack_0[128] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[128]/vcasc
+ bias_nstack
Xbias_nstack_0[129] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[129]/vcasc
+ bias_nstack
Xbias_nstack_0[130] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[130]/vcasc
+ bias_nstack
Xbias_nstack_0[131] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[131]/vcasc
+ bias_nstack
Xbias_nstack_0[132] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[132]/vcasc
+ bias_nstack
Xbias_nstack_0[133] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[133]/vcasc
+ bias_nstack
Xbias_nstack_0[134] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[134]/vcasc
+ bias_nstack
Xbias_nstack_0[135] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[135]/vcasc
+ bias_nstack
Xbias_nstack_0[136] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[136]/vcasc
+ bias_nstack
Xbias_nstack_0[137] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[137]/vcasc
+ bias_nstack
Xbias_nstack_0[138] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[138]/vcasc
+ bias_nstack
Xbias_nstack_0[139] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[139]/vcasc
+ bias_nstack
Xbias_nstack_0[140] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[140]/vcasc
+ bias_nstack
Xbias_nstack_0[141] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[141]/vcasc
+ bias_nstack
Xbias_nstack_0[142] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[142]/vcasc
+ bias_nstack
Xbias_nstack_0[143] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[143]/vcasc
+ bias_nstack
Xbias_nstack_0[144] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[144]/vcasc
+ bias_nstack
Xbias_nstack_0[145] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[145]/vcasc
+ bias_nstack
Xbias_nstack_0[146] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[146]/vcasc
+ bias_nstack
Xbias_nstack_0[147] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[147]/vcasc
+ bias_nstack
Xbias_nstack_0[148] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[148]/vcasc
+ bias_nstack
Xbias_nstack_0[149] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[149]/vcasc
+ bias_nstack
Xbias_nstack_0[150] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[150]/vcasc
+ bias_nstack
Xbias_nstack_0[151] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[151]/vcasc
+ bias_nstack
Xbias_nstack_0[152] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[152]/vcasc
+ bias_nstack
Xbias_nstack_0[153] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[153]/vcasc
+ bias_nstack
Xbias_nstack_0[154] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[154]/vcasc
+ bias_nstack
Xbias_nstack_0[155] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[155]/vcasc
+ bias_nstack
Xbias_nstack_0[156] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[156]/vcasc
+ bias_nstack
Xbias_nstack_0[157] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[157]/vcasc
+ bias_nstack
Xbias_nstack_0[158] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[158]/vcasc
+ bias_nstack
Xbias_nstack_0[159] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[159]/vcasc
+ bias_nstack
Xbias_nstack_0[160] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[160]/vcasc
+ bias_nstack
Xbias_nstack_0[161] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[161]/vcasc
+ bias_nstack
Xbias_nstack_0[162] snk_5000_0 ena_5000_0 bias_nstack_0[9]/nbias avss bias_nstack_0[162]/vcasc
+ bias_nstack
Xbias_nstack_0[163] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[163]/vcasc
+ bias_nstack
Xbias_nstack_0[164] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[164]/vcasc
+ bias_nstack
Xbias_nstack_0[165] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[165]/vcasc
+ bias_nstack
Xbias_nstack_0[166] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[166]/vcasc
+ bias_nstack
Xbias_nstack_0[167] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[167]/vcasc
+ bias_nstack
Xbias_nstack_0[168] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[168]/vcasc
+ bias_nstack
Xbias_nstack_0[169] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[169]/vcasc
+ bias_nstack
Xbias_nstack_0[170] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[170]/vcasc
+ bias_nstack
Xbias_nstack_0[171] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[171]/vcasc
+ bias_nstack
Xbias_nstack_0[172] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[172]/vcasc
+ bias_nstack
Xbias_nstack_0[173] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[173]/vcasc
+ bias_nstack
Xbias_nstack_0[174] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[174]/vcasc
+ bias_nstack
Xbias_nstack_0[175] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[175]/vcasc
+ bias_nstack
Xbias_nstack_0[176] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[176]/vcasc
+ bias_nstack
Xbias_nstack_0[177] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[177]/vcasc
+ bias_nstack
Xbias_nstack_0[178] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[178]/vcasc
+ bias_nstack
Xbias_nstack_0[179] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[179]/vcasc
+ bias_nstack
Xbias_nstack_0[180] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[180]/vcasc
+ bias_nstack
Xbias_nstack_0[181] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[181]/vcasc
+ bias_nstack
Xbias_nstack_0[182] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[182]/vcasc
+ bias_nstack
Xbias_nstack_0[183] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[183]/vcasc
+ bias_nstack
Xbias_nstack_0[184] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[184]/vcasc
+ bias_nstack
Xbias_nstack_0[185] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[185]/vcasc
+ bias_nstack
Xbias_nstack_0[186] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[186]/vcasc
+ bias_nstack
Xbias_nstack_0[187] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[187]/vcasc
+ bias_nstack
Xbias_nstack_0[188] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[188]/vcasc
+ bias_nstack
Xbias_nstack_0[189] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[189]/vcasc
+ bias_nstack
Xbias_nstack_0[190] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[190]/vcasc
+ bias_nstack
Xbias_nstack_0[191] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[191]/vcasc
+ bias_nstack
Xbias_nstack_0[192] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[192]/vcasc
+ bias_nstack
Xbias_nstack_0[193] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[193]/vcasc
+ bias_nstack
Xbias_nstack_0[194] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[194]/vcasc
+ bias_nstack
Xbias_nstack_0[195] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[195]/vcasc
+ bias_nstack
Xbias_nstack_0[196] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[196]/vcasc
+ bias_nstack
Xbias_nstack_0[197] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[197]/vcasc
+ bias_nstack
Xbias_nstack_0[198] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[198]/vcasc
+ bias_nstack
Xbias_nstack_0[199] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[199]/vcasc
+ bias_nstack
Xbias_nstack_0[200] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[200]/vcasc
+ bias_nstack
Xbias_nstack_0[201] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[201]/vcasc
+ bias_nstack
Xbias_nstack_0[202] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[202]/vcasc
+ bias_nstack
Xbias_nstack_0[203] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[203]/vcasc
+ bias_nstack
Xbias_nstack_0[204] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[204]/vcasc
+ bias_nstack
Xbias_nstack_0[205] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[205]/vcasc
+ bias_nstack
Xbias_nstack_0[206] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[206]/vcasc
+ bias_nstack
Xbias_nstack_0[207] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[207]/vcasc
+ bias_nstack
Xbias_nstack_0[208] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[208]/vcasc
+ bias_nstack
Xbias_nstack_0[209] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[209]/vcasc
+ bias_nstack
Xbias_nstack_0[210] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[210]/vcasc
+ bias_nstack
Xbias_nstack_0[211] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[211]/vcasc
+ bias_nstack
Xbias_nstack_0[212] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[212]/vcasc
+ bias_nstack
Xbias_nstack_0[213] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[213]/vcasc
+ bias_nstack
Xbias_nstack_0[214] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[214]/vcasc
+ bias_nstack
Xbias_nstack_0[215] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[215]/vcasc
+ bias_nstack
Xbias_nstack_0[216] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[216]/vcasc
+ bias_nstack
Xbias_nstack_0[217] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[217]/vcasc
+ bias_nstack
Xbias_nstack_0[218] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[218]/vcasc
+ bias_nstack
Xbias_nstack_0[219] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[219]/vcasc
+ bias_nstack
Xbias_nstack_0[220] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[220]/vcasc
+ bias_nstack
Xbias_nstack_0[221] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[221]/vcasc
+ bias_nstack
Xbias_nstack_0[222] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[222]/vcasc
+ bias_nstack
Xbias_nstack_0[223] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[223]/vcasc
+ bias_nstack
Xbias_nstack_0[224] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[224]/vcasc
+ bias_nstack
Xbias_nstack_0[225] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[225]/vcasc
+ bias_nstack
Xbias_nstack_0[226] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[226]/vcasc
+ bias_nstack
Xbias_nstack_0[227] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[227]/vcasc
+ bias_nstack
Xbias_nstack_0[228] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[228]/vcasc
+ bias_nstack
Xbias_nstack_0[229] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[229]/vcasc
+ bias_nstack
Xbias_nstack_0[230] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[230]/vcasc
+ bias_nstack
Xbias_nstack_0[231] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[231]/vcasc
+ bias_nstack
Xbias_nstack_0[232] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[232]/vcasc
+ bias_nstack
Xbias_nstack_0[233] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[233]/vcasc
+ bias_nstack
Xbias_nstack_0[234] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[234]/vcasc
+ bias_nstack
Xbias_nstack_0[235] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[235]/vcasc
+ bias_nstack
Xbias_nstack_0[236] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[236]/vcasc
+ bias_nstack
Xbias_nstack_0[237] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[237]/vcasc
+ bias_nstack
Xbias_nstack_0[238] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[238]/vcasc
+ bias_nstack
Xbias_nstack_0[239] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[239]/vcasc
+ bias_nstack
Xbias_nstack_0[240] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[240]/vcasc
+ bias_nstack
Xbias_nstack_0[241] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[241]/vcasc
+ bias_nstack
Xbias_nstack_0[242] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[242]/vcasc
+ bias_nstack
Xbias_nstack_0[243] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[243]/vcasc
+ bias_nstack
Xbias_nstack_0[244] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[244]/vcasc
+ bias_nstack
Xbias_nstack_0[245] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[245]/vcasc
+ bias_nstack
Xbias_nstack_0[246] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[246]/vcasc
+ bias_nstack
Xbias_nstack_0[247] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[247]/vcasc
+ bias_nstack
Xbias_nstack_0[248] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[248]/vcasc
+ bias_nstack
Xbias_nstack_0[249] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[249]/vcasc
+ bias_nstack
Xbias_nstack_0[250] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[250]/vcasc
+ bias_nstack
Xbias_nstack_0[251] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[251]/vcasc
+ bias_nstack
Xbias_nstack_0[252] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[252]/vcasc
+ bias_nstack
Xbias_nstack_0[253] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[253]/vcasc
+ bias_nstack
Xbias_nstack_0[254] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[254]/vcasc
+ bias_nstack
Xbias_nstack_0[255] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[255]/vcasc
+ bias_nstack
Xbias_nstack_0[256] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[256]/vcasc
+ bias_nstack
Xbias_nstack_0[257] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[257]/vcasc
+ bias_nstack
Xbias_nstack_0[258] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[258]/vcasc
+ bias_nstack
Xbias_nstack_0[259] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[259]/vcasc
+ bias_nstack
Xbias_nstack_0[260] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[260]/vcasc
+ bias_nstack
Xbias_nstack_0[261] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[261]/vcasc
+ bias_nstack
Xbias_nstack_0[262] snk_5000_1 ena_5000_1 bias_nstack_0[9]/nbias avss bias_nstack_0[262]/vcasc
+ bias_nstack
Xbias_nstack_0[263] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[263]/vcasc
+ bias_nstack
Xbias_nstack_0[264] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[264]/vcasc
+ bias_nstack
Xbias_nstack_0[265] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[265]/vcasc
+ bias_nstack
Xbias_nstack_0[266] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[266]/vcasc
+ bias_nstack
Xbias_nstack_0[267] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[267]/vcasc
+ bias_nstack
Xbias_nstack_0[268] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[268]/vcasc
+ bias_nstack
Xbias_nstack_0[269] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[269]/vcasc
+ bias_nstack
Xbias_nstack_0[270] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[270]/vcasc
+ bias_nstack
Xbias_nstack_0[271] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[271]/vcasc
+ bias_nstack
Xbias_nstack_0[272] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[272]/vcasc
+ bias_nstack
Xbias_nstack_0[273] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[273]/vcasc
+ bias_nstack
Xbias_nstack_0[274] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[274]/vcasc
+ bias_nstack
Xbias_nstack_0[275] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[275]/vcasc
+ bias_nstack
Xbias_nstack_0[276] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[276]/vcasc
+ bias_nstack
Xbias_nstack_0[277] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[277]/vcasc
+ bias_nstack
Xbias_nstack_0[278] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[278]/vcasc
+ bias_nstack
Xbias_nstack_0[279] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[279]/vcasc
+ bias_nstack
Xbias_nstack_0[280] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[280]/vcasc
+ bias_nstack
Xbias_nstack_0[281] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[281]/vcasc
+ bias_nstack
Xbias_nstack_0[282] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[282]/vcasc
+ bias_nstack
Xbias_nstack_0[283] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[283]/vcasc
+ bias_nstack
Xbias_nstack_0[284] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[284]/vcasc
+ bias_nstack
Xbias_nstack_0[285] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[285]/vcasc
+ bias_nstack
Xbias_nstack_0[286] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[286]/vcasc
+ bias_nstack
Xbias_nstack_0[287] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[287]/vcasc
+ bias_nstack
Xbias_nstack_0[288] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[288]/vcasc
+ bias_nstack
Xbias_nstack_0[289] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[289]/vcasc
+ bias_nstack
Xbias_nstack_0[290] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[290]/vcasc
+ bias_nstack
Xbias_nstack_0[291] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[291]/vcasc
+ bias_nstack
Xbias_nstack_0[292] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[292]/vcasc
+ bias_nstack
Xbias_nstack_0[293] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[293]/vcasc
+ bias_nstack
Xbias_nstack_0[294] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[294]/vcasc
+ bias_nstack
Xbias_nstack_0[295] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[295]/vcasc
+ bias_nstack
Xbias_nstack_0[296] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[296]/vcasc
+ bias_nstack
Xbias_nstack_0[297] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[297]/vcasc
+ bias_nstack
Xbias_nstack_0[298] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[298]/vcasc
+ bias_nstack
Xbias_nstack_0[299] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[299]/vcasc
+ bias_nstack
Xbias_nstack_0[300] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[300]/vcasc
+ bias_nstack
Xbias_nstack_0[301] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[301]/vcasc
+ bias_nstack
Xbias_nstack_0[302] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[302]/vcasc
+ bias_nstack
Xbias_nstack_0[303] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[303]/vcasc
+ bias_nstack
Xbias_nstack_0[304] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[304]/vcasc
+ bias_nstack
Xbias_nstack_0[305] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[305]/vcasc
+ bias_nstack
Xbias_nstack_0[306] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[306]/vcasc
+ bias_nstack
Xbias_nstack_0[307] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[307]/vcasc
+ bias_nstack
Xbias_nstack_0[308] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[308]/vcasc
+ bias_nstack
Xbias_nstack_0[309] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[309]/vcasc
+ bias_nstack
Xbias_nstack_0[310] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[310]/vcasc
+ bias_nstack
Xbias_nstack_0[311] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[311]/vcasc
+ bias_nstack
Xbias_nstack_0[312] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[312]/vcasc
+ bias_nstack
Xbias_nstack_0[313] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[313]/vcasc
+ bias_nstack
Xbias_nstack_0[314] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[314]/vcasc
+ bias_nstack
Xbias_nstack_0[315] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[315]/vcasc
+ bias_nstack
Xbias_nstack_0[316] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[316]/vcasc
+ bias_nstack
Xbias_nstack_0[317] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[317]/vcasc
+ bias_nstack
Xbias_nstack_0[318] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[318]/vcasc
+ bias_nstack
Xbias_nstack_0[319] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[319]/vcasc
+ bias_nstack
Xbias_nstack_0[320] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[320]/vcasc
+ bias_nstack
Xbias_nstack_0[321] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[321]/vcasc
+ bias_nstack
Xbias_nstack_0[322] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[322]/vcasc
+ bias_nstack
Xbias_nstack_0[323] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[323]/vcasc
+ bias_nstack
Xbias_nstack_0[324] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[324]/vcasc
+ bias_nstack
Xbias_nstack_0[325] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[325]/vcasc
+ bias_nstack
Xbias_nstack_0[326] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[326]/vcasc
+ bias_nstack
Xbias_nstack_0[327] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[327]/vcasc
+ bias_nstack
Xbias_nstack_0[328] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[328]/vcasc
+ bias_nstack
Xbias_nstack_0[329] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[329]/vcasc
+ bias_nstack
Xbias_nstack_0[330] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[330]/vcasc
+ bias_nstack
Xbias_nstack_0[331] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[331]/vcasc
+ bias_nstack
Xbias_nstack_0[332] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[332]/vcasc
+ bias_nstack
Xbias_nstack_0[333] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[333]/vcasc
+ bias_nstack
Xbias_nstack_0[334] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[334]/vcasc
+ bias_nstack
Xbias_nstack_0[335] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[335]/vcasc
+ bias_nstack
Xbias_nstack_0[336] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[336]/vcasc
+ bias_nstack
Xbias_nstack_0[337] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[337]/vcasc
+ bias_nstack
Xbias_nstack_0[338] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[338]/vcasc
+ bias_nstack
Xbias_nstack_0[339] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[339]/vcasc
+ bias_nstack
Xbias_nstack_0[340] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[340]/vcasc
+ bias_nstack
Xbias_nstack_0[341] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[341]/vcasc
+ bias_nstack
Xbias_nstack_0[342] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[342]/vcasc
+ bias_nstack
Xbias_nstack_0[343] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[343]/vcasc
+ bias_nstack
Xbias_nstack_0[344] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[344]/vcasc
+ bias_nstack
Xbias_nstack_0[345] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[345]/vcasc
+ bias_nstack
Xbias_nstack_0[346] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[346]/vcasc
+ bias_nstack
Xbias_nstack_0[347] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[347]/vcasc
+ bias_nstack
Xbias_nstack_0[348] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[348]/vcasc
+ bias_nstack
Xbias_nstack_0[349] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[349]/vcasc
+ bias_nstack
Xbias_nstack_0[350] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[350]/vcasc
+ bias_nstack
Xbias_nstack_0[351] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[351]/vcasc
+ bias_nstack
Xbias_nstack_0[352] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[352]/vcasc
+ bias_nstack
Xbias_nstack_0[353] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[353]/vcasc
+ bias_nstack
Xbias_nstack_0[354] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[354]/vcasc
+ bias_nstack
Xbias_nstack_0[355] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[355]/vcasc
+ bias_nstack
Xbias_nstack_0[356] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[356]/vcasc
+ bias_nstack
Xbias_nstack_0[357] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[357]/vcasc
+ bias_nstack
Xbias_nstack_0[358] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[358]/vcasc
+ bias_nstack
Xbias_nstack_0[359] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[359]/vcasc
+ bias_nstack
Xbias_nstack_0[360] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[360]/vcasc
+ bias_nstack
Xbias_nstack_0[361] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[361]/vcasc
+ bias_nstack
Xbias_nstack_0[362] snk_5000_2 ena_5000_2 bias_nstack_0[9]/nbias avss bias_nstack_0[362]/vcasc
+ bias_nstack
Xbias_nstack_0[363] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[363]/vcasc
+ bias_nstack
Xbias_nstack_0[364] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[364]/vcasc
+ bias_nstack
Xbias_nstack_0[365] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[365]/vcasc
+ bias_nstack
Xbias_nstack_0[366] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[366]/vcasc
+ bias_nstack
Xbias_nstack_0[367] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[367]/vcasc
+ bias_nstack
Xbias_nstack_0[368] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[368]/vcasc
+ bias_nstack
Xbias_nstack_0[369] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[369]/vcasc
+ bias_nstack
Xbias_nstack_0[370] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[370]/vcasc
+ bias_nstack
Xbias_nstack_0[371] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[371]/vcasc
+ bias_nstack
Xbias_nstack_0[372] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[372]/vcasc
+ bias_nstack
Xbias_nstack_0[373] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[373]/vcasc
+ bias_nstack
Xbias_nstack_0[374] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[374]/vcasc
+ bias_nstack
Xbias_nstack_0[375] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[375]/vcasc
+ bias_nstack
Xbias_nstack_0[376] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[376]/vcasc
+ bias_nstack
Xbias_nstack_0[377] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[377]/vcasc
+ bias_nstack
Xbias_nstack_0[378] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[378]/vcasc
+ bias_nstack
Xbias_nstack_0[379] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[379]/vcasc
+ bias_nstack
Xbias_nstack_0[380] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[380]/vcasc
+ bias_nstack
Xbias_nstack_0[381] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[381]/vcasc
+ bias_nstack
Xbias_nstack_0[382] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[382]/vcasc
+ bias_nstack
Xbias_nstack_0[383] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[383]/vcasc
+ bias_nstack
Xbias_nstack_0[384] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[384]/vcasc
+ bias_nstack
Xbias_nstack_0[385] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[385]/vcasc
+ bias_nstack
Xbias_nstack_0[386] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[386]/vcasc
+ bias_nstack
Xbias_nstack_0[387] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[387]/vcasc
+ bias_nstack
Xbias_nstack_0[388] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[388]/vcasc
+ bias_nstack
Xbias_nstack_0[389] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[389]/vcasc
+ bias_nstack
Xbias_nstack_0[390] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[390]/vcasc
+ bias_nstack
Xbias_nstack_0[391] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[391]/vcasc
+ bias_nstack
Xbias_nstack_0[392] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[392]/vcasc
+ bias_nstack
Xbias_nstack_0[393] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[393]/vcasc
+ bias_nstack
Xbias_nstack_0[394] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[394]/vcasc
+ bias_nstack
Xbias_nstack_0[395] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[395]/vcasc
+ bias_nstack
Xbias_nstack_0[396] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[396]/vcasc
+ bias_nstack
Xbias_nstack_0[397] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[397]/vcasc
+ bias_nstack
Xbias_nstack_0[398] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[398]/vcasc
+ bias_nstack
Xbias_nstack_0[399] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[399]/vcasc
+ bias_nstack
Xbias_nstack_0[400] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[400]/vcasc
+ bias_nstack
Xbias_nstack_0[401] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[401]/vcasc
+ bias_nstack
Xbias_nstack_0[402] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[402]/vcasc
+ bias_nstack
Xbias_nstack_0[403] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[403]/vcasc
+ bias_nstack
Xbias_nstack_0[404] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[404]/vcasc
+ bias_nstack
Xbias_nstack_0[405] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[405]/vcasc
+ bias_nstack
Xbias_nstack_0[406] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[406]/vcasc
+ bias_nstack
Xbias_nstack_0[407] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[407]/vcasc
+ bias_nstack
Xbias_nstack_0[408] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[408]/vcasc
+ bias_nstack
Xbias_nstack_0[409] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[409]/vcasc
+ bias_nstack
Xbias_nstack_0[410] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[410]/vcasc
+ bias_nstack
Xbias_nstack_0[411] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[411]/vcasc
+ bias_nstack
Xbias_nstack_0[412] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[412]/vcasc
+ bias_nstack
Xbias_nstack_0[413] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[413]/vcasc
+ bias_nstack
Xbias_nstack_0[414] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[414]/vcasc
+ bias_nstack
Xbias_nstack_0[415] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[415]/vcasc
+ bias_nstack
Xbias_nstack_0[416] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[416]/vcasc
+ bias_nstack
Xbias_nstack_0[417] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[417]/vcasc
+ bias_nstack
Xbias_nstack_0[418] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[418]/vcasc
+ bias_nstack
Xbias_nstack_0[419] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[419]/vcasc
+ bias_nstack
Xbias_nstack_0[420] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[420]/vcasc
+ bias_nstack
Xbias_nstack_0[421] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[421]/vcasc
+ bias_nstack
Xbias_nstack_0[422] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[422]/vcasc
+ bias_nstack
Xbias_nstack_0[423] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[423]/vcasc
+ bias_nstack
Xbias_nstack_0[424] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[424]/vcasc
+ bias_nstack
Xbias_nstack_0[425] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[425]/vcasc
+ bias_nstack
Xbias_nstack_0[426] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[426]/vcasc
+ bias_nstack
Xbias_nstack_0[427] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[427]/vcasc
+ bias_nstack
Xbias_nstack_0[428] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[428]/vcasc
+ bias_nstack
Xbias_nstack_0[429] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[429]/vcasc
+ bias_nstack
Xbias_nstack_0[430] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[430]/vcasc
+ bias_nstack
Xbias_nstack_0[431] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[431]/vcasc
+ bias_nstack
Xbias_nstack_0[432] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[432]/vcasc
+ bias_nstack
Xbias_nstack_0[433] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[433]/vcasc
+ bias_nstack
Xbias_nstack_0[434] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[434]/vcasc
+ bias_nstack
Xbias_nstack_0[435] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[435]/vcasc
+ bias_nstack
Xbias_nstack_0[436] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[436]/vcasc
+ bias_nstack
Xbias_nstack_0[437] snk_3700 ena_3700 bias_nstack_0[9]/nbias avss bias_nstack_0[437]/vcasc
+ bias_nstack
Xbias_nstack_0[438] snk_test1 ena_test1 bias_nstack_0[9]/nbias avss bias_nstack_0[438]/vcasc
+ bias_nstack
Xbias_nstack_0[439] snk_test1 ena_test1 bias_nstack_0[9]/nbias avss bias_nstack_0[439]/vcasc
+ bias_nstack
XXR2 m1_6353_1231# m1_11831_n5169# m1_2369_1231# m1_10005_1231# m1_9175_n5169# m1_4527_n5169#
+ m1_5855_n5169# m1_5357_1231# m1_10835_n5169# m1_10337_1231# m1_8179_n5169# m1_5025_1231#
+ m1_2037_1231# m1_5523_n5169# m1_12163_n5169# ref_in m1_8345_1231# m1_211_n5169#
+ m1_11333_1231# m1_6353_1231# m1_2369_1231# m1_7183_n5169# m1_11167_n5169# m1_12495_n5169#
+ m1_1207_n5169# m1_8013_1231# m1_11001_1231# m1_10171_n5169# m1_11499_n5169# m1_11333_1231#
+ m1_n121_n5169# m1_6851_n5169# m1_2701_1231# m1_4029_1231# m1_n287_1231# m1_8345_1231#
+ m1_5855_n5169# m1_2203_n5169# m1_10669_1231# m1_875_n5169# m1_6021_1231# m1_10503_n5169#
+ m1_3199_n5169# m1_4361_1231# m1_1373_1231# m1_45_1231# bias_pstack_0[9]/pcasc m1_12163_n5169#
+ m1_1871_n5169# m1_9009_1231# m1_9507_n5169# m1_6685_1231# m1_4195_n5169# m1_11001_1231#
+ m1_11167_n5169# m1_5025_1231# m1_8511_n5169# m1_12329_1231# m1_4693_1231# m1_2867_n5169#
+ m1_1705_1231# m1_1539_n5169# m1_9341_1231# m1_5191_n5169# m1_11665_1231# m1_6519_n5169#
+ m1_6685_1231# m1_10171_n5169# m1_3863_n5169# m1_2535_n5169# m1_2037_1231# m1_7515_n5169#
+ m1_8677_1231# m1_9175_n5169# m1_6851_n5169# m1_3531_n5169# m1_1705_1231# m1_9009_1231#
+ m1_11997_1231# m1_11831_n5169# m1_4859_n5169# m1_n453_n5169# m1_3697_1231# m1_1871_n5169#
+ m1_8677_1231# m1_709_1231# m1_8179_n5169# m1_11665_1231# m1_7349_1231# m1_4527_n5169#
+ m1_543_n5169# m1_10835_n5169# m1_5523_n5169# m1_4029_1231# m1_2867_n5169# m1_1041_1231#
+ m1_7183_n5169# m1_5689_1231# m1_9673_1231# m1_12495_n5169# m1_6187_n5169# m1_211_n5169#
+ avss m1_9839_n5169# m1_3697_1231# m1_709_1231# m1_7017_1231# m1_10005_1231# m1_3863_n5169#
+ m1_n121_n5169# m1_4361_1231# m1_1373_1231# m1_11499_n5169# m1_5689_1231# m1_9673_1231#
+ m1_1207_n5169# bias_nstack_0[61]/itail m1_4859_n5169# m1_8843_n5169# m1_875_n5169#
+ m1_n453_n5169# m1_7017_1231# m1_10503_n5169# m1_1041_1231# m1_2203_n5169# m1_3033_1231#
+ m1_7847_n5169# m1_9507_n5169# m1_2701_1231# m1_9341_1231# m1_6187_n5169# m1_n287_1231#
+ m1_8013_1231# m1_12329_1231# m1_543_n5169# m1_3199_n5169# m1_6021_1231# m1_3365_1231#
+ m1_1539_n5169# m1_377_1231# bias_pstack_0[9]/pcasc m1_8511_n5169# m1_10669_1231#
+ m1_11997_1231# m1_9839_n5169# m1_4195_n5169# m1_2535_n5169# m1_45_1231# m1_5191_n5169#
+ m1_7515_n5169# m1_5357_1231# m1_8843_n5169# m1_6519_n5169# m1_3033_1231# m1_4693_1231#
+ m1_377_1231# m1_7349_1231# m1_7847_n5169# m1_10337_1231# m1_3531_n5169# m1_3365_1231#
+ sky130_fd_pr__res_high_po_0p35_P35QVK
Xbias_pstack_0[0] avdd avss bias_pstack_0[9]/pcasc enb_test0 src_test0 bias_pstack_0[0]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[1] avdd avss bias_pstack_0[9]/pcasc enb_test0 src_test0 bias_pstack_0[1]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[2] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[2]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[3] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[3]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[4] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[4]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[5] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[5]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[6] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[6]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[7] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[7]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[8] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[8]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[9] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[9]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[10] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[10]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[11] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[11]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[12] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[12]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[13] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[13]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[14] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[14]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[15] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[15]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[16] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[16]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[17] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[17]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[18] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[18]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[19] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[19]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[20] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[20]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[21] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[21]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[22] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[22]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[23] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[23]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[24] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[24]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[25] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[25]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[26] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[26]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[27] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[27]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[28] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[28]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[29] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[29]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[30] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[30]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[31] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[31]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[32] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[32]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[33] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[33]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[34] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[34]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[35] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[35]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[36] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[36]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[37] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[37]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[38] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[38]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[39] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[39]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[40] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[40]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[41] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[41]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[42] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[42]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[43] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[43]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[44] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[44]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[45] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[45]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[46] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[46]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[47] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[47]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[48] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[48]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[49] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[49]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[50] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[50]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[51] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[51]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[52] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[52]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[53] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[53]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[54] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[54]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[55] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[55]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[56] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[56]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[57] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[57]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[58] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[58]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[59] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[59]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[60] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[60]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[61] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[61]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[62] avdd avss bias_pstack_0[9]/pcasc enb bias_pstack_0[62]/itail bias_pstack_0[9]/pbias
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[63] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[63]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[64] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[64]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[65] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[65]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[66] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[66]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[67] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[67]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[68] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[68]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[69] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[69]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[70] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[70]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[71] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[71]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[72] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[72]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[73] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[73]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[74] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[74]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[75] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[75]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[76] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[76]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[77] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[77]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[78] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[78]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[79] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[79]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[80] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[80]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[81] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[81]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[82] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[82]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[83] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[83]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[84] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[84]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[85] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[85]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[86] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[86]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[87] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[87]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[88] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[88]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[89] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[89]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[90] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[90]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[91] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[91]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[92] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[92]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[93] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[93]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[94] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[94]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[95] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[95]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[96] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[96]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[97] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[97]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[98] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[98]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[99] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[99]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[100] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[100]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[101] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[101]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[102] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[102]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[103] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[103]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[104] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[104]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[105] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[105]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[106] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[106]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[107] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[107]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[108] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[108]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[109] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[109]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[110] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[110]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[111] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[111]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[112] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[112]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[113] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[113]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[114] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[114]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[115] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[115]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[116] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[116]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[117] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[117]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[118] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[118]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[119] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[119]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[120] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[120]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[121] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[121]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[122] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[122]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[123] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[123]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[124] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[124]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[125] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[125]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[126] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[126]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[127] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[127]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[128] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[128]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[129] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[129]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[130] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[130]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[131] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[131]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[132] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[132]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[133] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[133]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[134] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[134]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[135] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[135]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[136] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[136]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[137] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[137]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[138] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[138]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[139] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[139]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[140] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[140]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[141] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[141]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[142] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[142]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[143] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[143]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[144] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[144]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[145] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[145]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[146] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[146]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[147] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[147]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[148] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[148]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[149] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[149]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[150] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[150]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[151] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[151]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[152] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[152]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[153] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[153]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[154] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[154]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[155] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[155]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[156] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[156]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[157] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[157]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[158] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[158]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[159] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[159]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[160] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[160]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[161] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[161]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[162] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[162]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[163] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[163]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[164] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[164]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[165] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[165]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[166] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[166]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[167] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[167]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[168] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[168]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[169] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[169]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[170] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[170]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[171] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[171]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[172] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[172]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[173] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[173]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[174] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[174]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[175] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[175]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[176] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[176]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[177] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[177]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[178] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[178]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[179] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[179]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[180] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[180]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[181] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[181]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[182] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[182]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[183] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[183]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[184] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[184]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[185] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[185]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[186] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[186]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[187] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[187]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[188] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[188]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[189] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[189]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[190] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[190]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[191] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[191]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[192] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[192]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[193] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[193]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[194] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[194]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[195] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[195]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[196] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[196]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[197] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[197]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[198] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[198]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[199] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[199]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[200] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[200]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[201] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[201]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[202] avdd avss bias_pstack_0[9]/pcasc enb_10000_0 src_10000_0 bias_pstack_0[202]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[203] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[203]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[204] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[204]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[205] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[205]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[206] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[206]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[207] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[207]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[208] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[208]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[209] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[209]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[210] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[210]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[211] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[211]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[212] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[212]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[213] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[213]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[214] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[214]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[215] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[215]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[216] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[216]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[217] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[217]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[218] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[218]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[219] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[219]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[220] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[220]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[221] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[221]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[222] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[222]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[223] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[223]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[224] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[224]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[225] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[225]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[226] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[226]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[227] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[227]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[228] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[228]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[229] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[229]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[230] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[230]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[231] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[231]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[232] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[232]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[233] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[233]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[234] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[234]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[235] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[235]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[236] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[236]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[237] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[237]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[238] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[238]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[239] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[239]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[240] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[240]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[241] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[241]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[242] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[242]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[243] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[243]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[244] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[244]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[245] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[245]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[246] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[246]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[247] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[247]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[248] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[248]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[249] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[249]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[250] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[250]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[251] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[251]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[252] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[252]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[253] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[253]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[254] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[254]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[255] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[255]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[256] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[256]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[257] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[257]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[258] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[258]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[259] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[259]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[260] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[260]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[261] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[261]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[262] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[262]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[263] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[263]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[264] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[264]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[265] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[265]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[266] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[266]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[267] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[267]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[268] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[268]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[269] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[269]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[270] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[270]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[271] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[271]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[272] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[272]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[273] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[273]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[274] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[274]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[275] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[275]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[276] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[276]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[277] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[277]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[278] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[278]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[279] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[279]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[280] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[280]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[281] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[281]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[282] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[282]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[283] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[283]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[284] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[284]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[285] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[285]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[286] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[286]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[287] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[287]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[288] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[288]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[289] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[289]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[290] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[290]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[291] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[291]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[292] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[292]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[293] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[293]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[294] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[294]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[295] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[295]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[296] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[296]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[297] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[297]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[298] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[298]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[299] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[299]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[300] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[300]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[301] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[301]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[302] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[302]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[303] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[303]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[304] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[304]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[305] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[305]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[306] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[306]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[307] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[307]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[308] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[308]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[309] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[309]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[310] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[310]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[311] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[311]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[312] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[312]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[313] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[313]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[314] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[314]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[315] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[315]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[316] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[316]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[317] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[317]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[318] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[318]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[319] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[319]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[320] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[320]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[321] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[321]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[322] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[322]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[323] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[323]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[324] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[324]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[325] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[325]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[326] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[326]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[327] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[327]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[328] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[328]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[329] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[329]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[330] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[330]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[331] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[331]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[332] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[332]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[333] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[333]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[334] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[334]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[335] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[335]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[336] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[336]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[337] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[337]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[338] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[338]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[339] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[339]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[340] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[340]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[341] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[341]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[342] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[342]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[343] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[343]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[344] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[344]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[345] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[345]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[346] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[346]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[347] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[347]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[348] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[348]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[349] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[349]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[350] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[350]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[351] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[351]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[352] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[352]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[353] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[353]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[354] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[354]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[355] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[355]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[356] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[356]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[357] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[357]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[358] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[358]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[359] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[359]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[360] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[360]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[361] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[361]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[362] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[362]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[363] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[363]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[364] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[364]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[365] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[365]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[366] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[366]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[367] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[367]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[368] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[368]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[369] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[369]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[370] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[370]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[371] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[371]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[372] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[372]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[373] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[373]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[374] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[374]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[375] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[375]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[376] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[376]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[377] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[377]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[378] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[378]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[379] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[379]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[380] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[380]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[381] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[381]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[382] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[382]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[383] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[383]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[384] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[384]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[385] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[385]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[386] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[386]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[387] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[387]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[388] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[388]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[389] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[389]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[390] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[390]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[391] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[391]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[392] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[392]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[393] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[393]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[394] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[394]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[395] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[395]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[396] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[396]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[397] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[397]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[398] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[398]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[399] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[399]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[400] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[400]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[401] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[401]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[402] avdd avss bias_pstack_0[9]/pcasc enb_10000_1 src_10000_1 bias_pstack_0[402]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[403] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[403]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[404] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[404]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[405] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[405]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[406] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[406]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[407] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[407]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[408] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[408]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[409] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[409]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[410] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[410]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[411] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[411]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[412] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[412]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[413] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[413]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[414] avdd avss bias_pstack_0[9]/pcasc enb_600 src_600 bias_pstack_0[414]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[415] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[415]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[416] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[416]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[417] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[417]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[418] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[418]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[419] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[419]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[420] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[420]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[421] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[421]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[422] avdd avss bias_pstack_0[9]/pcasc enb_400 src_400 bias_pstack_0[422]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[423] avdd avss bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[423]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[424] avdd avss bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[424]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[425] avdd avss bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[425]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[426] avdd avss bias_pstack_0[9]/pcasc enb_200_0 src_200_0 bias_pstack_0[426]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[427] avdd avss bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[427]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[428] avdd avss bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[428]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[429] avdd avss bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[429]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[430] avdd avss bias_pstack_0[9]/pcasc enb_200_1 src_200_1 bias_pstack_0[430]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[431] avdd avss bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[431]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[432] avdd avss bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[432]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[433] avdd avss bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[433]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[434] avdd avss bias_pstack_0[9]/pcasc enb_200_2 src_200_2 bias_pstack_0[434]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[435] avdd avss bias_pstack_0[9]/pcasc enb_100 src_100 bias_pstack_0[435]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[436] avdd avss bias_pstack_0[9]/pcasc enb_100 src_100 bias_pstack_0[436]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[437] avdd avss bias_pstack_0[9]/pcasc enb_50 src_50 bias_pstack_0[437]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[438] avdd avss bias_pstack_0[9]/pcasc enb_test1 src_test1 bias_pstack_0[438]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
Xbias_pstack_0[439] avdd avss bias_pstack_0[9]/pcasc enb_test1 src_test1 bias_pstack_0[439]/vcasc
+ bias_pstack_0[9]/pbias bias_pstack
.ends

