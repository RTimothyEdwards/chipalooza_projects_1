** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i
+ wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31] wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26]
+ wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23] wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16]
+ wbs_dat_i[15] wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7] wbs_dat_i[6]
+ wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31] wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28]
+ wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23] wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18]
+ wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15] wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8]
+ wbs_adr_i[7] wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o wbs_dat_o[31] wbs_dat_o[30]
+ wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24] wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20]
+ wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16] wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10]
+ wbs_dat_o[9] wbs_dat_o[8] wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121] la_data_in[120] la_data_in[119]
+ la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114] la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110]
+ la_data_in[109] la_data_in[108] la_data_in[107] la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101]
+ la_data_in[100] la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93] la_data_in[92]
+ la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86] la_data_in[85] la_data_in[84] la_data_in[83]
+ la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79] la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74]
+ la_data_in[73] la_data_in[72] la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58] la_data_in[57] la_data_in[56]
+ la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51] la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47]
+ la_data_in[46] la_data_in[45] la_data_in[44] la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38]
+ la_data_in[37] la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30] la_data_in[29]
+ la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23] la_data_in[22] la_data_in[21] la_data_in[20]
+ la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16] la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11]
+ la_data_in[10] la_data_in[9] la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123] la_data_out[122] la_data_out[121]
+ la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117] la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113]
+ la_data_out[112] la_data_out[111] la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98] la_data_out[97]
+ la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91] la_data_out[90] la_data_out[89] la_data_out[88]
+ la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84] la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79]
+ la_data_out[78] la_data_out[77] la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63] la_data_out[62] la_data_out[61]
+ la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56] la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52]
+ la_data_out[51] la_data_out[50] la_data_out[49] la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43]
+ la_data_out[42] la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35] la_data_out[34]
+ la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28] la_data_out[27] la_data_out[26] la_data_out[25]
+ la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21] la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16]
+ la_data_out[15] la_data_out[14] la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] la_oenb[127] la_oenb[126] la_oenb[125]
+ la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119] la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114]
+ la_oenb[113] la_oenb[112] la_oenb[111] la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94] la_oenb[93] la_oenb[92]
+ la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85] la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81]
+ la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76] la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70]
+ la_oenb[69] la_oenb[68] la_oenb[67] la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59]
+ la_oenb[58] la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49] la_oenb[48]
+ la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40] la_oenb[39] la_oenb[38] la_oenb[37]
+ la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31] la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26]
+ la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22] la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15]
+ la_oenb[14] la_oenb[13] la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4] la_oenb[3]
+ la_oenb[2] la_oenb[1] la_oenb[0] io_in[26] io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17]
+ io_in[16] io_in[15] io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4] io_in[3]
+ io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22] io_in_3v3[21] io_in_3v3[20] io_in_3v3[19]
+ io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14] io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9]
+ io_in_3v3[8] io_in_3v3[7] io_in_3v3[6] io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15] io_out[14] io_out[13]
+ io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5] io_out[4] io_out[3] io_out[2] io_out[1] io_out[0]
+ io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22] io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15]
+ io_oeb[14] io_oeb[13] io_oeb[12] io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13] gpio_analog[12] gpio_analog[11]
+ gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6] gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2]
+ gpio_analog[1] gpio_analog[0] gpio_noesd[17] gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11]
+ gpio_noesd[10] gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2] gpio_noesd[1]
+ gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5] io_analog[4] io_analog[3] io_analog[2]
+ io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1] io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_clock2
+ user_irq[2] user_irq[1] user_irq[0]
*.PININFO vdda1:B vdda2:B vssa1:B vssa2:B vccd1:B vccd2:B vssd1:B vssd2:B wb_clk_i:I wb_rst_i:I wbs_stb_i:I wbs_cyc_i:I wbs_we_i:I
*+ wbs_sel_i[3:0]:I wbs_dat_i[31:0]:I wbs_adr_i[31:0]:I wbs_ack_o:O wbs_dat_o[31:0]:O la_data_in[127:0]:I la_data_out[127:0]:O io_in[26:0]:I
*+ io_in_3v3[26:0]:I user_clock2:I io_out[26:0]:O io_oeb[26:0]:O gpio_analog[17:0]:B gpio_noesd[17:0]:B io_analog[10:0]:B io_clamp_high[2:0]:B
*+ io_clamp_low[2:0]:B user_irq[2:0]:O la_oenb[127:0]:I
x1 vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22] io_oeb[21] io_oeb[20] io_oeb[19]
+ io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12] io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6]
+ io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2] io_oeb[1] io_oeb[0] io_out[26] io_out[25] io_out[24] io_out[23] io_out[22] io_out[21] io_out[20]
+ io_out[19] io_out[18] io_out[17] io_out[16] io_out[15] io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7]
+ io_out[6] io_out[5] io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] gpio_noesd[17] gpio_noesd[16] gpio_noesd[15] gpio_noesd[14]
+ gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10] gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4]
+ gpio_noesd[3] gpio_noesd[2] gpio_noesd[1] gpio_noesd[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6] gpio_analog[5] gpio_analog[4]
+ gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124]
+ la_data_out[123] la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117] la_data_out[116]
+ la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111] la_data_out[110] la_data_out[109] la_data_out[108]
+ la_data_out[107] la_data_out[106] la_data_out[105] la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100]
+ la_data_out[99] la_data_out[98] la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84] la_data_out[83] la_data_out[82]
+ la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77] la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73]
+ la_data_out[72] la_data_out[71] la_data_out[70] la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64]
+ la_data_out[63] la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56] la_data_out[55]
+ la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49] la_data_out[48] la_data_out[47] la_data_out[46]
+ la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42] la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37]
+ la_data_out[36] la_data_out[35] la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21] la_data_out[20] la_data_out[19]
+ la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14] la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10]
+ la_data_out[9] la_data_out[8] la_data_out[7] la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1]
+ la_data_out[0] la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121] la_data_in[120]
+ la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114] la_data_in[113] la_data_in[112] la_data_in[111]
+ la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107] la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102]
+ la_data_in[101] la_data_in[100] la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86] la_data_in[85] la_data_in[84]
+ la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79] la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75]
+ la_data_in[74] la_data_in[73] la_data_in[72] la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66]
+ la_data_in[65] la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58] la_data_in[57]
+ la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51] la_data_in[50] la_data_in[49] la_data_in[48]
+ la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44] la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39]
+ la_data_in[38] la_data_in[37] la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23] la_data_in[22] la_data_in[21]
+ la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16] la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12]
+ la_data_in[11] la_data_in[10] la_data_in[9] la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2]
+ la_data_in[1] la_data_in[0] vssd2 vssd1 chipalooza_testchip1
.ends

* expanding   symbol:  chipalooza_testchip1.sym # of pins=15
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza_testchip1.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza_testchip1.sch
.subckt chipalooza_testchip1 vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22] io_oeb[21]
+ io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12] io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8]
+ io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2] io_oeb[1] io_oeb[0] io_out[26] io_out[25] io_out[24] io_out[23] io_out[22]
+ io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15] io_out[14] io_out[13] io_out[12] io_out[11] io_out[10]
+ io_out[9] io_out[8] io_out[7] io_out[6] io_out[5] io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] gpio_noesd[17] gpio_noesd[16]
+ gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10] gpio_noesd[9] gpio_noesd[8] gpio_noesd[7]
+ gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2] gpio_noesd[1] gpio_noesd[0] gpio_analog[17] gpio_analog[16]
+ gpio_analog[15] gpio_analog[14] gpio_analog[13] gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7]
+ gpio_analog[6] gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] io_analog[10] io_analog[9] io_analog[8]
+ io_analog[7] io_analog[6] io_analog[5] io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] la_data_out[127] la_data_out[126]
+ la_data_out[125] la_data_out[124] la_data_out[123] la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118]
+ la_data_out[117] la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111] la_data_out[110]
+ la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105] la_data_out[104] la_data_out[103] la_data_out[102]
+ la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98] la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93]
+ la_data_out[92] la_data_out[91] la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77] la_data_out[76] la_data_out[75]
+ la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70] la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66]
+ la_data_out[65] la_data_out[64] la_data_out[63] la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57]
+ la_data_out[56] la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49] la_data_out[48]
+ la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42] la_data_out[41] la_data_out[40] la_data_out[39]
+ la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35] la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30]
+ la_data_out[29] la_data_out[28] la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14] la_data_out[13] la_data_out[12]
+ la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7] la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3]
+ la_data_out[2] la_data_out[1] la_data_out[0] la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122]
+ la_data_in[121] la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114] la_data_in[113]
+ la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107] la_data_in[106] la_data_in[105] la_data_in[104]
+ la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100] la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95]
+ la_data_in[94] la_data_in[93] la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79] la_data_in[78] la_data_in[77]
+ la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72] la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68]
+ la_data_in[67] la_data_in[66] la_data_in[65] la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59]
+ la_data_in[58] la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51] la_data_in[50]
+ la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44] la_data_in[43] la_data_in[42] la_data_in[41]
+ la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37] la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32]
+ la_data_in[31] la_data_in[30] la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16] la_data_in[15] la_data_in[14]
+ la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9] la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4]
+ la_data_in[3] la_data_in[2] la_data_in[1] la_data_in[0] vssd2 vssd1
*.PININFO vdda1:I vssa1:I vccd2:I vdda2:I vssa2:I gpio_noesd[17:0]:B gpio_analog[17:0]:B la_data_out[127:0]:I io_out[26:0]:O
*+ la_data_in[127:0]:O io_oeb[26:0]:O io_analog[10:0]:B vssd2:I vssd1:I vccd1:I
x1 vdda1 gpio_analog[17] la_data_out[48] la_data_out[41] la_data_out[44] la_data_out[40] la_data_out[42] la_data_out[38]
+ la_data_out[46] la_data_out[47] la_data_out[49] la_data_out[45] la_data_out[39] la_data_out[43] src_200_0 src_10000_0 src_400 src_600 src_test1
+ src_200_1 src_100 src_10000_1 src_50 src_test0 src_200_2 la_data_out[78] la_data_out[125] la_data_out[84] la_data_out[82] la_data_out[81]
+ la_data_out[83] la_data_out[80] ibias_nc3 ibias_nc1 snk_5000_1 snk_test1 snk_3700 ibias_nc2 snk_test0 la_data_out[79] vssa1 bias_generator
x2 la_data_out[62] la_data_out[63] vssa2 vdda2 vdd_spare_3 power_stage
x3 la_data_out[60] la_data_out[61] vssa2 vdda2 io_analog[10] power_stage
x4 la_data_out[58] la_data_out[59] vssa2 vccd2 io_analog[9] power_stage
x5 la_data_out[56] la_data_out[57] vssa2 vdda2 io_analog[8] power_stage
x6 la_data_out[54] la_data_out[55] vssa2 vdda2 io_analog[7] power_stage
x7 la_data_out[52] la_data_out[53] vssa2 vdda2 io_analog[6] power_stage
x8 la_data_out[50] la_data_out[51] vssa2 vccd2 io_analog[5] power_stage
x9 la_data_out[65] la_data_out[64] vssa1 vdda1 io_analog[4] power_stage
x10 la_data_out[67] la_data_out[66] vssa1 vdda1 vdd_spare_2 power_stage
x11 la_data_out[69] la_data_out[68] vssa1 vdda1 io_analog[3] power_stage
x12 la_data_out[71] la_data_out[70] vssa1 vdda1 vdd_spare_1 power_stage
x13 la_data_out[73] la_data_out[72] vssa1 vdda1 io_analog[2] power_stage
x14 la_data_out[75] la_data_out[74] vssa1 vdda1 io_analog[1] power_stage
x15 la_data_out[77] la_data_out[76] vssa1 vdda1 io_analog[0] power_stage
X17 net4 gpio_analog[13] src_10000_1 vssd2 vssa2 io_analog[7] net2 net1 net3 lpopamp
x18 io_analog[0] vssa1 io_out[0] vccd1 net13 vssd1 io_out[1] vbgB la_data_out[112] la_data_out[113] la_data_out[111] net14 net15
+ la_data_out[107] la_data_out[106] la_data_out[108] net16 la_data_out[109] la_data_out[115] net17 la_data_out[114] la_data_in[117] io_out[5]
+ la_data_out[116] la_data_out[110] src_200_0 sky130_ajc_ip__brownout
x19 io_analog[1] vssa1 vccd1 vssd1 vbgB io_out[6] net18 la_data_out[105] la_data_out[104] la_data_out[103] la_data_out[102] net19
+ la_data_out[100] la_data_out[101] src_200_1 sky130_ajc_ip__overvoltage
x20 io_analog[2] net20 io_out[8] vssa1 vccd1 io_out[7] vssd1 io_out[3] vbgB io_out[2] la_data_out[96] la_data_out[97]
+ la_data_out[98] net21 la_data_out[94] io_out[4] net22 la_data_out[93] la_data_out[92] la_data_in[120] la_data_in[119] la_data_out[99]
+ la_data_out[95] src_200_2 sky130_ajc_ip__por
x21 vccd2 io_analog[8] vssa2 net6 io_out[17] net5 la_data_out[28] la_data_out[29] la_data_out[30] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[33] la_data_out[32] la_data_out[31] src_400 sky130_ak_ip__comparator
x22 io_analog[3] vssa1 vccd1 vssd1 src_50 la_data_out[86] la_data_out[85] io_out[12] gpio_noesd[3] gpio_noesd[4]
+ sky130_be_ip__lsxo
X23 gpio_analog[15] gpio_analog[14] la_data_out[19] la_data_out[20] io_out[23] io_analog[6] vccd2 vssa2 vssd2 src_10000_0 vssd2
+ sky130_ht_ip__hsxo_cpz1
x25 io_analog[10] gpio_noesd[7] src_100 net10 net9 vssa2 vccd2 vssd2 la_data_out[37] sky130_td_ip__opamp_hp
x26 io_analog[4] vccd1 la_data_out[91] la_data_out[87] src_600 la_data_out[88] io_out[13] vbgA la_data_out[89] la_data_out[90]
+ vssd1 vssa1 sky130_vbl_ip__overvoltage
x28 la_data_out[21] net1 net2 vccd2 vssd2 vdda2 lvl_shift_invert
x29 vssa2 la_data_out[22] net5 vdda2 net3 gpio_analog[12] vccd2 vssd2 analog_mux_sel1v8
x30 vssa2 la_data_out[23] net6 vdda2 net4 gpio_analog[11] vccd2 vssd2 analog_mux_sel1v8
x31 vccd2 vssd2 vssa2 la_data_out[17] gpio_analog[10] src_test1 vdda2 isolated_switch_ena1v8
x32 net8 io_analog[9] vssd2 vbgA la_data_out[35] net7 sky130_od_ip__tempsensor_ext_vp
x24 vssa2 la_data_out[34] net9 vdda2 net7 gpio_analog[9] vccd2 vssd2 analog_mux_sel1v8
x33 vssa2 la_data_out[36] net10 vdda2 net8 gpio_analog[8] vccd2 vssd2 analog_mux_sel1v8
x34 vccd1 vssd1 vssa1 la_data_out[124] gpio_analog[6] snk_test1 vdda1 isolated_switch_ena1v8
x35 vccd1 vssd1 vssa1 la_data_out[123] gpio_analog[5] snk_3700 vdda1 isolated_switch_ena1v8
x36 vssa1 la_data_out[122] vbgA vdda1 vbgB gpio_noesd[2] vccd1 vssd1 analog_mux_sel1v8
x37 vccd1 vssd1 vssa1 la_data_out[121] gpio_analog[1] snk_5000_1 vdda1 isolated_switch_ena1v8
x38 vccd1 vssd1 vssa1 la_data_out[118] gpio_analog[0] snk_test0 vdda1 isolated_switch_ena1v8
x16 io_analog[5] net12 vssd2 net11 la_data_out[9] la_data_out[8] la_data_out[10] la_data_out[7] la_data_out[11] la_data_out[6]
+ la_data_out[12] la_data_out[5] la_data_out[13] la_data_out[4] la_data_out[14] la_data_out[3] la_data_out[15] la_data_out[2] la_data_out[16]
+ la_data_out[1] bandgap
x39 io_analog[5] vssd2 net23 net11 bias_basis_current
x40 vssa2 la_data_out[18] net12 vdda2 src_test0 gpio_analog[16] vccd2 vssd2 analog_mux_sel1v8
R39 io_oeb[23] vssd2 0 m=1
R40 io_oeb[17] vssd2 0 m=1
R41 io_oeb[0] vssd1 0 m=1
R42 io_oeb[1] vssd1 0 m=1
R43 io_oeb[2] vssd1 0 m=1
R44 io_oeb[3] vssd1 0 m=1
R45 io_oeb[4] vssd1 0 m=1
R46 io_oeb[5] vssd1 0 m=1
R47 io_oeb[6] vssd1 0 m=1
R48 io_oeb[7] vssd1 0 m=1
R49 io_oeb[8] vssd1 0 m=1
R50 io_oeb[12] vssd1 0 m=1
R51 io_oeb[13] vssd1 0 m=1
.ends


* expanding   symbol:  bias_generator.sym # of pins=41
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/bias_generator.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/bias_generator.sch
.subckt bias_generator avdd ref_in enb enb_200_2 enb_400 enb_100 enb_200_1 enb_test1 enb_10000_1 enb_10000_0 enb_test0 enb_600
+ enb_50 enb_200_0 src_200_0 src_10000_0 src_400 src_600 src_test1 src_200_1 src_100 src_10000_1 src_50 src_test0 src_200_2 ena_test0
+ ena_2000 ena_test1 ena_5000_2 ena_5000_1 ena_3700 ena_5000_0 snk_5000_2 snk_2000 snk_5000_1 snk_test1 snk_3700 snk_5000_0 snk_test0 ena
+ avss
*.PININFO ref_in:I avss:B ena:I enb:I avdd:B enb_test0:I ena_test0:I src_test0:B snk_test0:B ena_test1:I snk_test1:B enb_test1:I
*+ src_test1:B enb_10000_0:I src_10000_0:B ena_5000_0:I snk_5000_0:B enb_10000_1:I src_10000_1:B ena_5000_1:I snk_5000_1:B ena_5000_2:I
*+ snk_5000_2:B enb_600:I src_600:B enb_400:I src_400:B enb_200_0:I src_200_0:B enb_200_1:I src_200_1:B enb_200_2:I src_200_2:B enb_100:I
*+ src_100:B enb_50:I src_50:B ena_3700:I snk_3700:B ena_2000:I snk_2000:B
x2[19] net1 ena nbias nbias avss bias_nstack
x2[18] net1 ena nbias nbias avss bias_nstack
x2[17] net1 ena nbias nbias avss bias_nstack
x2[16] net1 ena nbias nbias avss bias_nstack
x2[15] net1 ena nbias nbias avss bias_nstack
x2[14] net1 ena nbias nbias avss bias_nstack
x2[13] net1 ena nbias nbias avss bias_nstack
x2[12] net1 ena nbias nbias avss bias_nstack
x2[11] net1 ena nbias nbias avss bias_nstack
x2[10] net1 ena nbias nbias avss bias_nstack
x2[9] net1 ena nbias nbias avss bias_nstack
x2[8] net1 ena nbias nbias avss bias_nstack
x2[7] net1 ena nbias nbias avss bias_nstack
x2[6] net1 ena nbias nbias avss bias_nstack
x2[5] net1 ena nbias nbias avss bias_nstack
x2[4] net1 ena nbias nbias avss bias_nstack
x2[3] net1 ena nbias nbias avss bias_nstack
x2[2] net1 ena nbias nbias avss bias_nstack
x2[1] net1 ena nbias nbias avss bias_nstack
x2[0] net1 ena nbias nbias avss bias_nstack
XR3 net1 pcasc avss sky130_fd_pr__res_high_po_0p35 L=900 mult=1 m=1
XR4 pcasc ref_in avss sky130_fd_pr__res_high_po_0p35 L=1500 mult=1 m=1
x4 net2 ena net3 nbias avss bias_nstack
x2 avdd pbias pcasc pbias enb avss net2 bias_pstack
x13[1] avdd pbias pcasc net4[1] enb_test0 avss src_test0 bias_pstack
x13[0] avdd pbias pcasc net4[0] enb_test0 avss src_test0 bias_pstack
x17[1] snk_test0 ena_test0 net5[1] nbias avss bias_nstack
x17[0] snk_test0 ena_test0 net5[0] nbias avss bias_nstack
x18[1] snk_test1 ena_test1 net6[1] nbias avss bias_nstack
x18[0] snk_test1 ena_test1 net6[0] nbias avss bias_nstack
x16[1] avdd pbias pcasc net7[1] enb_test1 avss src_test1 bias_pstack
x16[0] avdd pbias pcasc net7[0] enb_test1 avss src_test1 bias_pstack
x8[199] avdd pbias pcasc net8[199] enb_10000_0 avss src_10000_0 bias_pstack
x8[198] avdd pbias pcasc net8[198] enb_10000_0 avss src_10000_0 bias_pstack
x8[197] avdd pbias pcasc net8[197] enb_10000_0 avss src_10000_0 bias_pstack
x8[196] avdd pbias pcasc net8[196] enb_10000_0 avss src_10000_0 bias_pstack
x8[195] avdd pbias pcasc net8[195] enb_10000_0 avss src_10000_0 bias_pstack
x8[194] avdd pbias pcasc net8[194] enb_10000_0 avss src_10000_0 bias_pstack
x8[193] avdd pbias pcasc net8[193] enb_10000_0 avss src_10000_0 bias_pstack
x8[192] avdd pbias pcasc net8[192] enb_10000_0 avss src_10000_0 bias_pstack
x8[191] avdd pbias pcasc net8[191] enb_10000_0 avss src_10000_0 bias_pstack
x8[190] avdd pbias pcasc net8[190] enb_10000_0 avss src_10000_0 bias_pstack
x8[189] avdd pbias pcasc net8[189] enb_10000_0 avss src_10000_0 bias_pstack
x8[188] avdd pbias pcasc net8[188] enb_10000_0 avss src_10000_0 bias_pstack
x8[187] avdd pbias pcasc net8[187] enb_10000_0 avss src_10000_0 bias_pstack
x8[186] avdd pbias pcasc net8[186] enb_10000_0 avss src_10000_0 bias_pstack
x8[185] avdd pbias pcasc net8[185] enb_10000_0 avss src_10000_0 bias_pstack
x8[184] avdd pbias pcasc net8[184] enb_10000_0 avss src_10000_0 bias_pstack
x8[183] avdd pbias pcasc net8[183] enb_10000_0 avss src_10000_0 bias_pstack
x8[182] avdd pbias pcasc net8[182] enb_10000_0 avss src_10000_0 bias_pstack
x8[181] avdd pbias pcasc net8[181] enb_10000_0 avss src_10000_0 bias_pstack
x8[180] avdd pbias pcasc net8[180] enb_10000_0 avss src_10000_0 bias_pstack
x8[179] avdd pbias pcasc net8[179] enb_10000_0 avss src_10000_0 bias_pstack
x8[178] avdd pbias pcasc net8[178] enb_10000_0 avss src_10000_0 bias_pstack
x8[177] avdd pbias pcasc net8[177] enb_10000_0 avss src_10000_0 bias_pstack
x8[176] avdd pbias pcasc net8[176] enb_10000_0 avss src_10000_0 bias_pstack
x8[175] avdd pbias pcasc net8[175] enb_10000_0 avss src_10000_0 bias_pstack
x8[174] avdd pbias pcasc net8[174] enb_10000_0 avss src_10000_0 bias_pstack
x8[173] avdd pbias pcasc net8[173] enb_10000_0 avss src_10000_0 bias_pstack
x8[172] avdd pbias pcasc net8[172] enb_10000_0 avss src_10000_0 bias_pstack
x8[171] avdd pbias pcasc net8[171] enb_10000_0 avss src_10000_0 bias_pstack
x8[170] avdd pbias pcasc net8[170] enb_10000_0 avss src_10000_0 bias_pstack
x8[169] avdd pbias pcasc net8[169] enb_10000_0 avss src_10000_0 bias_pstack
x8[168] avdd pbias pcasc net8[168] enb_10000_0 avss src_10000_0 bias_pstack
x8[167] avdd pbias pcasc net8[167] enb_10000_0 avss src_10000_0 bias_pstack
x8[166] avdd pbias pcasc net8[166] enb_10000_0 avss src_10000_0 bias_pstack
x8[165] avdd pbias pcasc net8[165] enb_10000_0 avss src_10000_0 bias_pstack
x8[164] avdd pbias pcasc net8[164] enb_10000_0 avss src_10000_0 bias_pstack
x8[163] avdd pbias pcasc net8[163] enb_10000_0 avss src_10000_0 bias_pstack
x8[162] avdd pbias pcasc net8[162] enb_10000_0 avss src_10000_0 bias_pstack
x8[161] avdd pbias pcasc net8[161] enb_10000_0 avss src_10000_0 bias_pstack
x8[160] avdd pbias pcasc net8[160] enb_10000_0 avss src_10000_0 bias_pstack
x8[159] avdd pbias pcasc net8[159] enb_10000_0 avss src_10000_0 bias_pstack
x8[158] avdd pbias pcasc net8[158] enb_10000_0 avss src_10000_0 bias_pstack
x8[157] avdd pbias pcasc net8[157] enb_10000_0 avss src_10000_0 bias_pstack
x8[156] avdd pbias pcasc net8[156] enb_10000_0 avss src_10000_0 bias_pstack
x8[155] avdd pbias pcasc net8[155] enb_10000_0 avss src_10000_0 bias_pstack
x8[154] avdd pbias pcasc net8[154] enb_10000_0 avss src_10000_0 bias_pstack
x8[153] avdd pbias pcasc net8[153] enb_10000_0 avss src_10000_0 bias_pstack
x8[152] avdd pbias pcasc net8[152] enb_10000_0 avss src_10000_0 bias_pstack
x8[151] avdd pbias pcasc net8[151] enb_10000_0 avss src_10000_0 bias_pstack
x8[150] avdd pbias pcasc net8[150] enb_10000_0 avss src_10000_0 bias_pstack
x8[149] avdd pbias pcasc net8[149] enb_10000_0 avss src_10000_0 bias_pstack
x8[148] avdd pbias pcasc net8[148] enb_10000_0 avss src_10000_0 bias_pstack
x8[147] avdd pbias pcasc net8[147] enb_10000_0 avss src_10000_0 bias_pstack
x8[146] avdd pbias pcasc net8[146] enb_10000_0 avss src_10000_0 bias_pstack
x8[145] avdd pbias pcasc net8[145] enb_10000_0 avss src_10000_0 bias_pstack
x8[144] avdd pbias pcasc net8[144] enb_10000_0 avss src_10000_0 bias_pstack
x8[143] avdd pbias pcasc net8[143] enb_10000_0 avss src_10000_0 bias_pstack
x8[142] avdd pbias pcasc net8[142] enb_10000_0 avss src_10000_0 bias_pstack
x8[141] avdd pbias pcasc net8[141] enb_10000_0 avss src_10000_0 bias_pstack
x8[140] avdd pbias pcasc net8[140] enb_10000_0 avss src_10000_0 bias_pstack
x8[139] avdd pbias pcasc net8[139] enb_10000_0 avss src_10000_0 bias_pstack
x8[138] avdd pbias pcasc net8[138] enb_10000_0 avss src_10000_0 bias_pstack
x8[137] avdd pbias pcasc net8[137] enb_10000_0 avss src_10000_0 bias_pstack
x8[136] avdd pbias pcasc net8[136] enb_10000_0 avss src_10000_0 bias_pstack
x8[135] avdd pbias pcasc net8[135] enb_10000_0 avss src_10000_0 bias_pstack
x8[134] avdd pbias pcasc net8[134] enb_10000_0 avss src_10000_0 bias_pstack
x8[133] avdd pbias pcasc net8[133] enb_10000_0 avss src_10000_0 bias_pstack
x8[132] avdd pbias pcasc net8[132] enb_10000_0 avss src_10000_0 bias_pstack
x8[131] avdd pbias pcasc net8[131] enb_10000_0 avss src_10000_0 bias_pstack
x8[130] avdd pbias pcasc net8[130] enb_10000_0 avss src_10000_0 bias_pstack
x8[129] avdd pbias pcasc net8[129] enb_10000_0 avss src_10000_0 bias_pstack
x8[128] avdd pbias pcasc net8[128] enb_10000_0 avss src_10000_0 bias_pstack
x8[127] avdd pbias pcasc net8[127] enb_10000_0 avss src_10000_0 bias_pstack
x8[126] avdd pbias pcasc net8[126] enb_10000_0 avss src_10000_0 bias_pstack
x8[125] avdd pbias pcasc net8[125] enb_10000_0 avss src_10000_0 bias_pstack
x8[124] avdd pbias pcasc net8[124] enb_10000_0 avss src_10000_0 bias_pstack
x8[123] avdd pbias pcasc net8[123] enb_10000_0 avss src_10000_0 bias_pstack
x8[122] avdd pbias pcasc net8[122] enb_10000_0 avss src_10000_0 bias_pstack
x8[121] avdd pbias pcasc net8[121] enb_10000_0 avss src_10000_0 bias_pstack
x8[120] avdd pbias pcasc net8[120] enb_10000_0 avss src_10000_0 bias_pstack
x8[119] avdd pbias pcasc net8[119] enb_10000_0 avss src_10000_0 bias_pstack
x8[118] avdd pbias pcasc net8[118] enb_10000_0 avss src_10000_0 bias_pstack
x8[117] avdd pbias pcasc net8[117] enb_10000_0 avss src_10000_0 bias_pstack
x8[116] avdd pbias pcasc net8[116] enb_10000_0 avss src_10000_0 bias_pstack
x8[115] avdd pbias pcasc net8[115] enb_10000_0 avss src_10000_0 bias_pstack
x8[114] avdd pbias pcasc net8[114] enb_10000_0 avss src_10000_0 bias_pstack
x8[113] avdd pbias pcasc net8[113] enb_10000_0 avss src_10000_0 bias_pstack
x8[112] avdd pbias pcasc net8[112] enb_10000_0 avss src_10000_0 bias_pstack
x8[111] avdd pbias pcasc net8[111] enb_10000_0 avss src_10000_0 bias_pstack
x8[110] avdd pbias pcasc net8[110] enb_10000_0 avss src_10000_0 bias_pstack
x8[109] avdd pbias pcasc net8[109] enb_10000_0 avss src_10000_0 bias_pstack
x8[108] avdd pbias pcasc net8[108] enb_10000_0 avss src_10000_0 bias_pstack
x8[107] avdd pbias pcasc net8[107] enb_10000_0 avss src_10000_0 bias_pstack
x8[106] avdd pbias pcasc net8[106] enb_10000_0 avss src_10000_0 bias_pstack
x8[105] avdd pbias pcasc net8[105] enb_10000_0 avss src_10000_0 bias_pstack
x8[104] avdd pbias pcasc net8[104] enb_10000_0 avss src_10000_0 bias_pstack
x8[103] avdd pbias pcasc net8[103] enb_10000_0 avss src_10000_0 bias_pstack
x8[102] avdd pbias pcasc net8[102] enb_10000_0 avss src_10000_0 bias_pstack
x8[101] avdd pbias pcasc net8[101] enb_10000_0 avss src_10000_0 bias_pstack
x8[100] avdd pbias pcasc net8[100] enb_10000_0 avss src_10000_0 bias_pstack
x8[99] avdd pbias pcasc net8[99] enb_10000_0 avss src_10000_0 bias_pstack
x8[98] avdd pbias pcasc net8[98] enb_10000_0 avss src_10000_0 bias_pstack
x8[97] avdd pbias pcasc net8[97] enb_10000_0 avss src_10000_0 bias_pstack
x8[96] avdd pbias pcasc net8[96] enb_10000_0 avss src_10000_0 bias_pstack
x8[95] avdd pbias pcasc net8[95] enb_10000_0 avss src_10000_0 bias_pstack
x8[94] avdd pbias pcasc net8[94] enb_10000_0 avss src_10000_0 bias_pstack
x8[93] avdd pbias pcasc net8[93] enb_10000_0 avss src_10000_0 bias_pstack
x8[92] avdd pbias pcasc net8[92] enb_10000_0 avss src_10000_0 bias_pstack
x8[91] avdd pbias pcasc net8[91] enb_10000_0 avss src_10000_0 bias_pstack
x8[90] avdd pbias pcasc net8[90] enb_10000_0 avss src_10000_0 bias_pstack
x8[89] avdd pbias pcasc net8[89] enb_10000_0 avss src_10000_0 bias_pstack
x8[88] avdd pbias pcasc net8[88] enb_10000_0 avss src_10000_0 bias_pstack
x8[87] avdd pbias pcasc net8[87] enb_10000_0 avss src_10000_0 bias_pstack
x8[86] avdd pbias pcasc net8[86] enb_10000_0 avss src_10000_0 bias_pstack
x8[85] avdd pbias pcasc net8[85] enb_10000_0 avss src_10000_0 bias_pstack
x8[84] avdd pbias pcasc net8[84] enb_10000_0 avss src_10000_0 bias_pstack
x8[83] avdd pbias pcasc net8[83] enb_10000_0 avss src_10000_0 bias_pstack
x8[82] avdd pbias pcasc net8[82] enb_10000_0 avss src_10000_0 bias_pstack
x8[81] avdd pbias pcasc net8[81] enb_10000_0 avss src_10000_0 bias_pstack
x8[80] avdd pbias pcasc net8[80] enb_10000_0 avss src_10000_0 bias_pstack
x8[79] avdd pbias pcasc net8[79] enb_10000_0 avss src_10000_0 bias_pstack
x8[78] avdd pbias pcasc net8[78] enb_10000_0 avss src_10000_0 bias_pstack
x8[77] avdd pbias pcasc net8[77] enb_10000_0 avss src_10000_0 bias_pstack
x8[76] avdd pbias pcasc net8[76] enb_10000_0 avss src_10000_0 bias_pstack
x8[75] avdd pbias pcasc net8[75] enb_10000_0 avss src_10000_0 bias_pstack
x8[74] avdd pbias pcasc net8[74] enb_10000_0 avss src_10000_0 bias_pstack
x8[73] avdd pbias pcasc net8[73] enb_10000_0 avss src_10000_0 bias_pstack
x8[72] avdd pbias pcasc net8[72] enb_10000_0 avss src_10000_0 bias_pstack
x8[71] avdd pbias pcasc net8[71] enb_10000_0 avss src_10000_0 bias_pstack
x8[70] avdd pbias pcasc net8[70] enb_10000_0 avss src_10000_0 bias_pstack
x8[69] avdd pbias pcasc net8[69] enb_10000_0 avss src_10000_0 bias_pstack
x8[68] avdd pbias pcasc net8[68] enb_10000_0 avss src_10000_0 bias_pstack
x8[67] avdd pbias pcasc net8[67] enb_10000_0 avss src_10000_0 bias_pstack
x8[66] avdd pbias pcasc net8[66] enb_10000_0 avss src_10000_0 bias_pstack
x8[65] avdd pbias pcasc net8[65] enb_10000_0 avss src_10000_0 bias_pstack
x8[64] avdd pbias pcasc net8[64] enb_10000_0 avss src_10000_0 bias_pstack
x8[63] avdd pbias pcasc net8[63] enb_10000_0 avss src_10000_0 bias_pstack
x8[62] avdd pbias pcasc net8[62] enb_10000_0 avss src_10000_0 bias_pstack
x8[61] avdd pbias pcasc net8[61] enb_10000_0 avss src_10000_0 bias_pstack
x8[60] avdd pbias pcasc net8[60] enb_10000_0 avss src_10000_0 bias_pstack
x8[59] avdd pbias pcasc net8[59] enb_10000_0 avss src_10000_0 bias_pstack
x8[58] avdd pbias pcasc net8[58] enb_10000_0 avss src_10000_0 bias_pstack
x8[57] avdd pbias pcasc net8[57] enb_10000_0 avss src_10000_0 bias_pstack
x8[56] avdd pbias pcasc net8[56] enb_10000_0 avss src_10000_0 bias_pstack
x8[55] avdd pbias pcasc net8[55] enb_10000_0 avss src_10000_0 bias_pstack
x8[54] avdd pbias pcasc net8[54] enb_10000_0 avss src_10000_0 bias_pstack
x8[53] avdd pbias pcasc net8[53] enb_10000_0 avss src_10000_0 bias_pstack
x8[52] avdd pbias pcasc net8[52] enb_10000_0 avss src_10000_0 bias_pstack
x8[51] avdd pbias pcasc net8[51] enb_10000_0 avss src_10000_0 bias_pstack
x8[50] avdd pbias pcasc net8[50] enb_10000_0 avss src_10000_0 bias_pstack
x8[49] avdd pbias pcasc net8[49] enb_10000_0 avss src_10000_0 bias_pstack
x8[48] avdd pbias pcasc net8[48] enb_10000_0 avss src_10000_0 bias_pstack
x8[47] avdd pbias pcasc net8[47] enb_10000_0 avss src_10000_0 bias_pstack
x8[46] avdd pbias pcasc net8[46] enb_10000_0 avss src_10000_0 bias_pstack
x8[45] avdd pbias pcasc net8[45] enb_10000_0 avss src_10000_0 bias_pstack
x8[44] avdd pbias pcasc net8[44] enb_10000_0 avss src_10000_0 bias_pstack
x8[43] avdd pbias pcasc net8[43] enb_10000_0 avss src_10000_0 bias_pstack
x8[42] avdd pbias pcasc net8[42] enb_10000_0 avss src_10000_0 bias_pstack
x8[41] avdd pbias pcasc net8[41] enb_10000_0 avss src_10000_0 bias_pstack
x8[40] avdd pbias pcasc net8[40] enb_10000_0 avss src_10000_0 bias_pstack
x8[39] avdd pbias pcasc net8[39] enb_10000_0 avss src_10000_0 bias_pstack
x8[38] avdd pbias pcasc net8[38] enb_10000_0 avss src_10000_0 bias_pstack
x8[37] avdd pbias pcasc net8[37] enb_10000_0 avss src_10000_0 bias_pstack
x8[36] avdd pbias pcasc net8[36] enb_10000_0 avss src_10000_0 bias_pstack
x8[35] avdd pbias pcasc net8[35] enb_10000_0 avss src_10000_0 bias_pstack
x8[34] avdd pbias pcasc net8[34] enb_10000_0 avss src_10000_0 bias_pstack
x8[33] avdd pbias pcasc net8[33] enb_10000_0 avss src_10000_0 bias_pstack
x8[32] avdd pbias pcasc net8[32] enb_10000_0 avss src_10000_0 bias_pstack
x8[31] avdd pbias pcasc net8[31] enb_10000_0 avss src_10000_0 bias_pstack
x8[30] avdd pbias pcasc net8[30] enb_10000_0 avss src_10000_0 bias_pstack
x8[29] avdd pbias pcasc net8[29] enb_10000_0 avss src_10000_0 bias_pstack
x8[28] avdd pbias pcasc net8[28] enb_10000_0 avss src_10000_0 bias_pstack
x8[27] avdd pbias pcasc net8[27] enb_10000_0 avss src_10000_0 bias_pstack
x8[26] avdd pbias pcasc net8[26] enb_10000_0 avss src_10000_0 bias_pstack
x8[25] avdd pbias pcasc net8[25] enb_10000_0 avss src_10000_0 bias_pstack
x8[24] avdd pbias pcasc net8[24] enb_10000_0 avss src_10000_0 bias_pstack
x8[23] avdd pbias pcasc net8[23] enb_10000_0 avss src_10000_0 bias_pstack
x8[22] avdd pbias pcasc net8[22] enb_10000_0 avss src_10000_0 bias_pstack
x8[21] avdd pbias pcasc net8[21] enb_10000_0 avss src_10000_0 bias_pstack
x8[20] avdd pbias pcasc net8[20] enb_10000_0 avss src_10000_0 bias_pstack
x8[19] avdd pbias pcasc net8[19] enb_10000_0 avss src_10000_0 bias_pstack
x8[18] avdd pbias pcasc net8[18] enb_10000_0 avss src_10000_0 bias_pstack
x8[17] avdd pbias pcasc net8[17] enb_10000_0 avss src_10000_0 bias_pstack
x8[16] avdd pbias pcasc net8[16] enb_10000_0 avss src_10000_0 bias_pstack
x8[15] avdd pbias pcasc net8[15] enb_10000_0 avss src_10000_0 bias_pstack
x8[14] avdd pbias pcasc net8[14] enb_10000_0 avss src_10000_0 bias_pstack
x8[13] avdd pbias pcasc net8[13] enb_10000_0 avss src_10000_0 bias_pstack
x8[12] avdd pbias pcasc net8[12] enb_10000_0 avss src_10000_0 bias_pstack
x8[11] avdd pbias pcasc net8[11] enb_10000_0 avss src_10000_0 bias_pstack
x8[10] avdd pbias pcasc net8[10] enb_10000_0 avss src_10000_0 bias_pstack
x8[9] avdd pbias pcasc net8[9] enb_10000_0 avss src_10000_0 bias_pstack
x8[8] avdd pbias pcasc net8[8] enb_10000_0 avss src_10000_0 bias_pstack
x8[7] avdd pbias pcasc net8[7] enb_10000_0 avss src_10000_0 bias_pstack
x8[6] avdd pbias pcasc net8[6] enb_10000_0 avss src_10000_0 bias_pstack
x8[5] avdd pbias pcasc net8[5] enb_10000_0 avss src_10000_0 bias_pstack
x8[4] avdd pbias pcasc net8[4] enb_10000_0 avss src_10000_0 bias_pstack
x8[3] avdd pbias pcasc net8[3] enb_10000_0 avss src_10000_0 bias_pstack
x8[2] avdd pbias pcasc net8[2] enb_10000_0 avss src_10000_0 bias_pstack
x8[1] avdd pbias pcasc net8[1] enb_10000_0 avss src_10000_0 bias_pstack
x8[0] avdd pbias pcasc net8[0] enb_10000_0 avss src_10000_0 bias_pstack
x9[99] snk_5000_0 ena_5000_0 net9[99] nbias avss bias_nstack
x9[98] snk_5000_0 ena_5000_0 net9[98] nbias avss bias_nstack
x9[97] snk_5000_0 ena_5000_0 net9[97] nbias avss bias_nstack
x9[96] snk_5000_0 ena_5000_0 net9[96] nbias avss bias_nstack
x9[95] snk_5000_0 ena_5000_0 net9[95] nbias avss bias_nstack
x9[94] snk_5000_0 ena_5000_0 net9[94] nbias avss bias_nstack
x9[93] snk_5000_0 ena_5000_0 net9[93] nbias avss bias_nstack
x9[92] snk_5000_0 ena_5000_0 net9[92] nbias avss bias_nstack
x9[91] snk_5000_0 ena_5000_0 net9[91] nbias avss bias_nstack
x9[90] snk_5000_0 ena_5000_0 net9[90] nbias avss bias_nstack
x9[89] snk_5000_0 ena_5000_0 net9[89] nbias avss bias_nstack
x9[88] snk_5000_0 ena_5000_0 net9[88] nbias avss bias_nstack
x9[87] snk_5000_0 ena_5000_0 net9[87] nbias avss bias_nstack
x9[86] snk_5000_0 ena_5000_0 net9[86] nbias avss bias_nstack
x9[85] snk_5000_0 ena_5000_0 net9[85] nbias avss bias_nstack
x9[84] snk_5000_0 ena_5000_0 net9[84] nbias avss bias_nstack
x9[83] snk_5000_0 ena_5000_0 net9[83] nbias avss bias_nstack
x9[82] snk_5000_0 ena_5000_0 net9[82] nbias avss bias_nstack
x9[81] snk_5000_0 ena_5000_0 net9[81] nbias avss bias_nstack
x9[80] snk_5000_0 ena_5000_0 net9[80] nbias avss bias_nstack
x9[79] snk_5000_0 ena_5000_0 net9[79] nbias avss bias_nstack
x9[78] snk_5000_0 ena_5000_0 net9[78] nbias avss bias_nstack
x9[77] snk_5000_0 ena_5000_0 net9[77] nbias avss bias_nstack
x9[76] snk_5000_0 ena_5000_0 net9[76] nbias avss bias_nstack
x9[75] snk_5000_0 ena_5000_0 net9[75] nbias avss bias_nstack
x9[74] snk_5000_0 ena_5000_0 net9[74] nbias avss bias_nstack
x9[73] snk_5000_0 ena_5000_0 net9[73] nbias avss bias_nstack
x9[72] snk_5000_0 ena_5000_0 net9[72] nbias avss bias_nstack
x9[71] snk_5000_0 ena_5000_0 net9[71] nbias avss bias_nstack
x9[70] snk_5000_0 ena_5000_0 net9[70] nbias avss bias_nstack
x9[69] snk_5000_0 ena_5000_0 net9[69] nbias avss bias_nstack
x9[68] snk_5000_0 ena_5000_0 net9[68] nbias avss bias_nstack
x9[67] snk_5000_0 ena_5000_0 net9[67] nbias avss bias_nstack
x9[66] snk_5000_0 ena_5000_0 net9[66] nbias avss bias_nstack
x9[65] snk_5000_0 ena_5000_0 net9[65] nbias avss bias_nstack
x9[64] snk_5000_0 ena_5000_0 net9[64] nbias avss bias_nstack
x9[63] snk_5000_0 ena_5000_0 net9[63] nbias avss bias_nstack
x9[62] snk_5000_0 ena_5000_0 net9[62] nbias avss bias_nstack
x9[61] snk_5000_0 ena_5000_0 net9[61] nbias avss bias_nstack
x9[60] snk_5000_0 ena_5000_0 net9[60] nbias avss bias_nstack
x9[59] snk_5000_0 ena_5000_0 net9[59] nbias avss bias_nstack
x9[58] snk_5000_0 ena_5000_0 net9[58] nbias avss bias_nstack
x9[57] snk_5000_0 ena_5000_0 net9[57] nbias avss bias_nstack
x9[56] snk_5000_0 ena_5000_0 net9[56] nbias avss bias_nstack
x9[55] snk_5000_0 ena_5000_0 net9[55] nbias avss bias_nstack
x9[54] snk_5000_0 ena_5000_0 net9[54] nbias avss bias_nstack
x9[53] snk_5000_0 ena_5000_0 net9[53] nbias avss bias_nstack
x9[52] snk_5000_0 ena_5000_0 net9[52] nbias avss bias_nstack
x9[51] snk_5000_0 ena_5000_0 net9[51] nbias avss bias_nstack
x9[50] snk_5000_0 ena_5000_0 net9[50] nbias avss bias_nstack
x9[49] snk_5000_0 ena_5000_0 net9[49] nbias avss bias_nstack
x9[48] snk_5000_0 ena_5000_0 net9[48] nbias avss bias_nstack
x9[47] snk_5000_0 ena_5000_0 net9[47] nbias avss bias_nstack
x9[46] snk_5000_0 ena_5000_0 net9[46] nbias avss bias_nstack
x9[45] snk_5000_0 ena_5000_0 net9[45] nbias avss bias_nstack
x9[44] snk_5000_0 ena_5000_0 net9[44] nbias avss bias_nstack
x9[43] snk_5000_0 ena_5000_0 net9[43] nbias avss bias_nstack
x9[42] snk_5000_0 ena_5000_0 net9[42] nbias avss bias_nstack
x9[41] snk_5000_0 ena_5000_0 net9[41] nbias avss bias_nstack
x9[40] snk_5000_0 ena_5000_0 net9[40] nbias avss bias_nstack
x9[39] snk_5000_0 ena_5000_0 net9[39] nbias avss bias_nstack
x9[38] snk_5000_0 ena_5000_0 net9[38] nbias avss bias_nstack
x9[37] snk_5000_0 ena_5000_0 net9[37] nbias avss bias_nstack
x9[36] snk_5000_0 ena_5000_0 net9[36] nbias avss bias_nstack
x9[35] snk_5000_0 ena_5000_0 net9[35] nbias avss bias_nstack
x9[34] snk_5000_0 ena_5000_0 net9[34] nbias avss bias_nstack
x9[33] snk_5000_0 ena_5000_0 net9[33] nbias avss bias_nstack
x9[32] snk_5000_0 ena_5000_0 net9[32] nbias avss bias_nstack
x9[31] snk_5000_0 ena_5000_0 net9[31] nbias avss bias_nstack
x9[30] snk_5000_0 ena_5000_0 net9[30] nbias avss bias_nstack
x9[29] snk_5000_0 ena_5000_0 net9[29] nbias avss bias_nstack
x9[28] snk_5000_0 ena_5000_0 net9[28] nbias avss bias_nstack
x9[27] snk_5000_0 ena_5000_0 net9[27] nbias avss bias_nstack
x9[26] snk_5000_0 ena_5000_0 net9[26] nbias avss bias_nstack
x9[25] snk_5000_0 ena_5000_0 net9[25] nbias avss bias_nstack
x9[24] snk_5000_0 ena_5000_0 net9[24] nbias avss bias_nstack
x9[23] snk_5000_0 ena_5000_0 net9[23] nbias avss bias_nstack
x9[22] snk_5000_0 ena_5000_0 net9[22] nbias avss bias_nstack
x9[21] snk_5000_0 ena_5000_0 net9[21] nbias avss bias_nstack
x9[20] snk_5000_0 ena_5000_0 net9[20] nbias avss bias_nstack
x9[19] snk_5000_0 ena_5000_0 net9[19] nbias avss bias_nstack
x9[18] snk_5000_0 ena_5000_0 net9[18] nbias avss bias_nstack
x9[17] snk_5000_0 ena_5000_0 net9[17] nbias avss bias_nstack
x9[16] snk_5000_0 ena_5000_0 net9[16] nbias avss bias_nstack
x9[15] snk_5000_0 ena_5000_0 net9[15] nbias avss bias_nstack
x9[14] snk_5000_0 ena_5000_0 net9[14] nbias avss bias_nstack
x9[13] snk_5000_0 ena_5000_0 net9[13] nbias avss bias_nstack
x9[12] snk_5000_0 ena_5000_0 net9[12] nbias avss bias_nstack
x9[11] snk_5000_0 ena_5000_0 net9[11] nbias avss bias_nstack
x9[10] snk_5000_0 ena_5000_0 net9[10] nbias avss bias_nstack
x9[9] snk_5000_0 ena_5000_0 net9[9] nbias avss bias_nstack
x9[8] snk_5000_0 ena_5000_0 net9[8] nbias avss bias_nstack
x9[7] snk_5000_0 ena_5000_0 net9[7] nbias avss bias_nstack
x9[6] snk_5000_0 ena_5000_0 net9[6] nbias avss bias_nstack
x9[5] snk_5000_0 ena_5000_0 net9[5] nbias avss bias_nstack
x9[4] snk_5000_0 ena_5000_0 net9[4] nbias avss bias_nstack
x9[3] snk_5000_0 ena_5000_0 net9[3] nbias avss bias_nstack
x9[2] snk_5000_0 ena_5000_0 net9[2] nbias avss bias_nstack
x9[1] snk_5000_0 ena_5000_0 net9[1] nbias avss bias_nstack
x9[0] snk_5000_0 ena_5000_0 net9[0] nbias avss bias_nstack
x10[199] avdd pbias pcasc net10[199] enb_10000_1 avss src_10000_1 bias_pstack
x10[198] avdd pbias pcasc net10[198] enb_10000_1 avss src_10000_1 bias_pstack
x10[197] avdd pbias pcasc net10[197] enb_10000_1 avss src_10000_1 bias_pstack
x10[196] avdd pbias pcasc net10[196] enb_10000_1 avss src_10000_1 bias_pstack
x10[195] avdd pbias pcasc net10[195] enb_10000_1 avss src_10000_1 bias_pstack
x10[194] avdd pbias pcasc net10[194] enb_10000_1 avss src_10000_1 bias_pstack
x10[193] avdd pbias pcasc net10[193] enb_10000_1 avss src_10000_1 bias_pstack
x10[192] avdd pbias pcasc net10[192] enb_10000_1 avss src_10000_1 bias_pstack
x10[191] avdd pbias pcasc net10[191] enb_10000_1 avss src_10000_1 bias_pstack
x10[190] avdd pbias pcasc net10[190] enb_10000_1 avss src_10000_1 bias_pstack
x10[189] avdd pbias pcasc net10[189] enb_10000_1 avss src_10000_1 bias_pstack
x10[188] avdd pbias pcasc net10[188] enb_10000_1 avss src_10000_1 bias_pstack
x10[187] avdd pbias pcasc net10[187] enb_10000_1 avss src_10000_1 bias_pstack
x10[186] avdd pbias pcasc net10[186] enb_10000_1 avss src_10000_1 bias_pstack
x10[185] avdd pbias pcasc net10[185] enb_10000_1 avss src_10000_1 bias_pstack
x10[184] avdd pbias pcasc net10[184] enb_10000_1 avss src_10000_1 bias_pstack
x10[183] avdd pbias pcasc net10[183] enb_10000_1 avss src_10000_1 bias_pstack
x10[182] avdd pbias pcasc net10[182] enb_10000_1 avss src_10000_1 bias_pstack
x10[181] avdd pbias pcasc net10[181] enb_10000_1 avss src_10000_1 bias_pstack
x10[180] avdd pbias pcasc net10[180] enb_10000_1 avss src_10000_1 bias_pstack
x10[179] avdd pbias pcasc net10[179] enb_10000_1 avss src_10000_1 bias_pstack
x10[178] avdd pbias pcasc net10[178] enb_10000_1 avss src_10000_1 bias_pstack
x10[177] avdd pbias pcasc net10[177] enb_10000_1 avss src_10000_1 bias_pstack
x10[176] avdd pbias pcasc net10[176] enb_10000_1 avss src_10000_1 bias_pstack
x10[175] avdd pbias pcasc net10[175] enb_10000_1 avss src_10000_1 bias_pstack
x10[174] avdd pbias pcasc net10[174] enb_10000_1 avss src_10000_1 bias_pstack
x10[173] avdd pbias pcasc net10[173] enb_10000_1 avss src_10000_1 bias_pstack
x10[172] avdd pbias pcasc net10[172] enb_10000_1 avss src_10000_1 bias_pstack
x10[171] avdd pbias pcasc net10[171] enb_10000_1 avss src_10000_1 bias_pstack
x10[170] avdd pbias pcasc net10[170] enb_10000_1 avss src_10000_1 bias_pstack
x10[169] avdd pbias pcasc net10[169] enb_10000_1 avss src_10000_1 bias_pstack
x10[168] avdd pbias pcasc net10[168] enb_10000_1 avss src_10000_1 bias_pstack
x10[167] avdd pbias pcasc net10[167] enb_10000_1 avss src_10000_1 bias_pstack
x10[166] avdd pbias pcasc net10[166] enb_10000_1 avss src_10000_1 bias_pstack
x10[165] avdd pbias pcasc net10[165] enb_10000_1 avss src_10000_1 bias_pstack
x10[164] avdd pbias pcasc net10[164] enb_10000_1 avss src_10000_1 bias_pstack
x10[163] avdd pbias pcasc net10[163] enb_10000_1 avss src_10000_1 bias_pstack
x10[162] avdd pbias pcasc net10[162] enb_10000_1 avss src_10000_1 bias_pstack
x10[161] avdd pbias pcasc net10[161] enb_10000_1 avss src_10000_1 bias_pstack
x10[160] avdd pbias pcasc net10[160] enb_10000_1 avss src_10000_1 bias_pstack
x10[159] avdd pbias pcasc net10[159] enb_10000_1 avss src_10000_1 bias_pstack
x10[158] avdd pbias pcasc net10[158] enb_10000_1 avss src_10000_1 bias_pstack
x10[157] avdd pbias pcasc net10[157] enb_10000_1 avss src_10000_1 bias_pstack
x10[156] avdd pbias pcasc net10[156] enb_10000_1 avss src_10000_1 bias_pstack
x10[155] avdd pbias pcasc net10[155] enb_10000_1 avss src_10000_1 bias_pstack
x10[154] avdd pbias pcasc net10[154] enb_10000_1 avss src_10000_1 bias_pstack
x10[153] avdd pbias pcasc net10[153] enb_10000_1 avss src_10000_1 bias_pstack
x10[152] avdd pbias pcasc net10[152] enb_10000_1 avss src_10000_1 bias_pstack
x10[151] avdd pbias pcasc net10[151] enb_10000_1 avss src_10000_1 bias_pstack
x10[150] avdd pbias pcasc net10[150] enb_10000_1 avss src_10000_1 bias_pstack
x10[149] avdd pbias pcasc net10[149] enb_10000_1 avss src_10000_1 bias_pstack
x10[148] avdd pbias pcasc net10[148] enb_10000_1 avss src_10000_1 bias_pstack
x10[147] avdd pbias pcasc net10[147] enb_10000_1 avss src_10000_1 bias_pstack
x10[146] avdd pbias pcasc net10[146] enb_10000_1 avss src_10000_1 bias_pstack
x10[145] avdd pbias pcasc net10[145] enb_10000_1 avss src_10000_1 bias_pstack
x10[144] avdd pbias pcasc net10[144] enb_10000_1 avss src_10000_1 bias_pstack
x10[143] avdd pbias pcasc net10[143] enb_10000_1 avss src_10000_1 bias_pstack
x10[142] avdd pbias pcasc net10[142] enb_10000_1 avss src_10000_1 bias_pstack
x10[141] avdd pbias pcasc net10[141] enb_10000_1 avss src_10000_1 bias_pstack
x10[140] avdd pbias pcasc net10[140] enb_10000_1 avss src_10000_1 bias_pstack
x10[139] avdd pbias pcasc net10[139] enb_10000_1 avss src_10000_1 bias_pstack
x10[138] avdd pbias pcasc net10[138] enb_10000_1 avss src_10000_1 bias_pstack
x10[137] avdd pbias pcasc net10[137] enb_10000_1 avss src_10000_1 bias_pstack
x10[136] avdd pbias pcasc net10[136] enb_10000_1 avss src_10000_1 bias_pstack
x10[135] avdd pbias pcasc net10[135] enb_10000_1 avss src_10000_1 bias_pstack
x10[134] avdd pbias pcasc net10[134] enb_10000_1 avss src_10000_1 bias_pstack
x10[133] avdd pbias pcasc net10[133] enb_10000_1 avss src_10000_1 bias_pstack
x10[132] avdd pbias pcasc net10[132] enb_10000_1 avss src_10000_1 bias_pstack
x10[131] avdd pbias pcasc net10[131] enb_10000_1 avss src_10000_1 bias_pstack
x10[130] avdd pbias pcasc net10[130] enb_10000_1 avss src_10000_1 bias_pstack
x10[129] avdd pbias pcasc net10[129] enb_10000_1 avss src_10000_1 bias_pstack
x10[128] avdd pbias pcasc net10[128] enb_10000_1 avss src_10000_1 bias_pstack
x10[127] avdd pbias pcasc net10[127] enb_10000_1 avss src_10000_1 bias_pstack
x10[126] avdd pbias pcasc net10[126] enb_10000_1 avss src_10000_1 bias_pstack
x10[125] avdd pbias pcasc net10[125] enb_10000_1 avss src_10000_1 bias_pstack
x10[124] avdd pbias pcasc net10[124] enb_10000_1 avss src_10000_1 bias_pstack
x10[123] avdd pbias pcasc net10[123] enb_10000_1 avss src_10000_1 bias_pstack
x10[122] avdd pbias pcasc net10[122] enb_10000_1 avss src_10000_1 bias_pstack
x10[121] avdd pbias pcasc net10[121] enb_10000_1 avss src_10000_1 bias_pstack
x10[120] avdd pbias pcasc net10[120] enb_10000_1 avss src_10000_1 bias_pstack
x10[119] avdd pbias pcasc net10[119] enb_10000_1 avss src_10000_1 bias_pstack
x10[118] avdd pbias pcasc net10[118] enb_10000_1 avss src_10000_1 bias_pstack
x10[117] avdd pbias pcasc net10[117] enb_10000_1 avss src_10000_1 bias_pstack
x10[116] avdd pbias pcasc net10[116] enb_10000_1 avss src_10000_1 bias_pstack
x10[115] avdd pbias pcasc net10[115] enb_10000_1 avss src_10000_1 bias_pstack
x10[114] avdd pbias pcasc net10[114] enb_10000_1 avss src_10000_1 bias_pstack
x10[113] avdd pbias pcasc net10[113] enb_10000_1 avss src_10000_1 bias_pstack
x10[112] avdd pbias pcasc net10[112] enb_10000_1 avss src_10000_1 bias_pstack
x10[111] avdd pbias pcasc net10[111] enb_10000_1 avss src_10000_1 bias_pstack
x10[110] avdd pbias pcasc net10[110] enb_10000_1 avss src_10000_1 bias_pstack
x10[109] avdd pbias pcasc net10[109] enb_10000_1 avss src_10000_1 bias_pstack
x10[108] avdd pbias pcasc net10[108] enb_10000_1 avss src_10000_1 bias_pstack
x10[107] avdd pbias pcasc net10[107] enb_10000_1 avss src_10000_1 bias_pstack
x10[106] avdd pbias pcasc net10[106] enb_10000_1 avss src_10000_1 bias_pstack
x10[105] avdd pbias pcasc net10[105] enb_10000_1 avss src_10000_1 bias_pstack
x10[104] avdd pbias pcasc net10[104] enb_10000_1 avss src_10000_1 bias_pstack
x10[103] avdd pbias pcasc net10[103] enb_10000_1 avss src_10000_1 bias_pstack
x10[102] avdd pbias pcasc net10[102] enb_10000_1 avss src_10000_1 bias_pstack
x10[101] avdd pbias pcasc net10[101] enb_10000_1 avss src_10000_1 bias_pstack
x10[100] avdd pbias pcasc net10[100] enb_10000_1 avss src_10000_1 bias_pstack
x10[99] avdd pbias pcasc net10[99] enb_10000_1 avss src_10000_1 bias_pstack
x10[98] avdd pbias pcasc net10[98] enb_10000_1 avss src_10000_1 bias_pstack
x10[97] avdd pbias pcasc net10[97] enb_10000_1 avss src_10000_1 bias_pstack
x10[96] avdd pbias pcasc net10[96] enb_10000_1 avss src_10000_1 bias_pstack
x10[95] avdd pbias pcasc net10[95] enb_10000_1 avss src_10000_1 bias_pstack
x10[94] avdd pbias pcasc net10[94] enb_10000_1 avss src_10000_1 bias_pstack
x10[93] avdd pbias pcasc net10[93] enb_10000_1 avss src_10000_1 bias_pstack
x10[92] avdd pbias pcasc net10[92] enb_10000_1 avss src_10000_1 bias_pstack
x10[91] avdd pbias pcasc net10[91] enb_10000_1 avss src_10000_1 bias_pstack
x10[90] avdd pbias pcasc net10[90] enb_10000_1 avss src_10000_1 bias_pstack
x10[89] avdd pbias pcasc net10[89] enb_10000_1 avss src_10000_1 bias_pstack
x10[88] avdd pbias pcasc net10[88] enb_10000_1 avss src_10000_1 bias_pstack
x10[87] avdd pbias pcasc net10[87] enb_10000_1 avss src_10000_1 bias_pstack
x10[86] avdd pbias pcasc net10[86] enb_10000_1 avss src_10000_1 bias_pstack
x10[85] avdd pbias pcasc net10[85] enb_10000_1 avss src_10000_1 bias_pstack
x10[84] avdd pbias pcasc net10[84] enb_10000_1 avss src_10000_1 bias_pstack
x10[83] avdd pbias pcasc net10[83] enb_10000_1 avss src_10000_1 bias_pstack
x10[82] avdd pbias pcasc net10[82] enb_10000_1 avss src_10000_1 bias_pstack
x10[81] avdd pbias pcasc net10[81] enb_10000_1 avss src_10000_1 bias_pstack
x10[80] avdd pbias pcasc net10[80] enb_10000_1 avss src_10000_1 bias_pstack
x10[79] avdd pbias pcasc net10[79] enb_10000_1 avss src_10000_1 bias_pstack
x10[78] avdd pbias pcasc net10[78] enb_10000_1 avss src_10000_1 bias_pstack
x10[77] avdd pbias pcasc net10[77] enb_10000_1 avss src_10000_1 bias_pstack
x10[76] avdd pbias pcasc net10[76] enb_10000_1 avss src_10000_1 bias_pstack
x10[75] avdd pbias pcasc net10[75] enb_10000_1 avss src_10000_1 bias_pstack
x10[74] avdd pbias pcasc net10[74] enb_10000_1 avss src_10000_1 bias_pstack
x10[73] avdd pbias pcasc net10[73] enb_10000_1 avss src_10000_1 bias_pstack
x10[72] avdd pbias pcasc net10[72] enb_10000_1 avss src_10000_1 bias_pstack
x10[71] avdd pbias pcasc net10[71] enb_10000_1 avss src_10000_1 bias_pstack
x10[70] avdd pbias pcasc net10[70] enb_10000_1 avss src_10000_1 bias_pstack
x10[69] avdd pbias pcasc net10[69] enb_10000_1 avss src_10000_1 bias_pstack
x10[68] avdd pbias pcasc net10[68] enb_10000_1 avss src_10000_1 bias_pstack
x10[67] avdd pbias pcasc net10[67] enb_10000_1 avss src_10000_1 bias_pstack
x10[66] avdd pbias pcasc net10[66] enb_10000_1 avss src_10000_1 bias_pstack
x10[65] avdd pbias pcasc net10[65] enb_10000_1 avss src_10000_1 bias_pstack
x10[64] avdd pbias pcasc net10[64] enb_10000_1 avss src_10000_1 bias_pstack
x10[63] avdd pbias pcasc net10[63] enb_10000_1 avss src_10000_1 bias_pstack
x10[62] avdd pbias pcasc net10[62] enb_10000_1 avss src_10000_1 bias_pstack
x10[61] avdd pbias pcasc net10[61] enb_10000_1 avss src_10000_1 bias_pstack
x10[60] avdd pbias pcasc net10[60] enb_10000_1 avss src_10000_1 bias_pstack
x10[59] avdd pbias pcasc net10[59] enb_10000_1 avss src_10000_1 bias_pstack
x10[58] avdd pbias pcasc net10[58] enb_10000_1 avss src_10000_1 bias_pstack
x10[57] avdd pbias pcasc net10[57] enb_10000_1 avss src_10000_1 bias_pstack
x10[56] avdd pbias pcasc net10[56] enb_10000_1 avss src_10000_1 bias_pstack
x10[55] avdd pbias pcasc net10[55] enb_10000_1 avss src_10000_1 bias_pstack
x10[54] avdd pbias pcasc net10[54] enb_10000_1 avss src_10000_1 bias_pstack
x10[53] avdd pbias pcasc net10[53] enb_10000_1 avss src_10000_1 bias_pstack
x10[52] avdd pbias pcasc net10[52] enb_10000_1 avss src_10000_1 bias_pstack
x10[51] avdd pbias pcasc net10[51] enb_10000_1 avss src_10000_1 bias_pstack
x10[50] avdd pbias pcasc net10[50] enb_10000_1 avss src_10000_1 bias_pstack
x10[49] avdd pbias pcasc net10[49] enb_10000_1 avss src_10000_1 bias_pstack
x10[48] avdd pbias pcasc net10[48] enb_10000_1 avss src_10000_1 bias_pstack
x10[47] avdd pbias pcasc net10[47] enb_10000_1 avss src_10000_1 bias_pstack
x10[46] avdd pbias pcasc net10[46] enb_10000_1 avss src_10000_1 bias_pstack
x10[45] avdd pbias pcasc net10[45] enb_10000_1 avss src_10000_1 bias_pstack
x10[44] avdd pbias pcasc net10[44] enb_10000_1 avss src_10000_1 bias_pstack
x10[43] avdd pbias pcasc net10[43] enb_10000_1 avss src_10000_1 bias_pstack
x10[42] avdd pbias pcasc net10[42] enb_10000_1 avss src_10000_1 bias_pstack
x10[41] avdd pbias pcasc net10[41] enb_10000_1 avss src_10000_1 bias_pstack
x10[40] avdd pbias pcasc net10[40] enb_10000_1 avss src_10000_1 bias_pstack
x10[39] avdd pbias pcasc net10[39] enb_10000_1 avss src_10000_1 bias_pstack
x10[38] avdd pbias pcasc net10[38] enb_10000_1 avss src_10000_1 bias_pstack
x10[37] avdd pbias pcasc net10[37] enb_10000_1 avss src_10000_1 bias_pstack
x10[36] avdd pbias pcasc net10[36] enb_10000_1 avss src_10000_1 bias_pstack
x10[35] avdd pbias pcasc net10[35] enb_10000_1 avss src_10000_1 bias_pstack
x10[34] avdd pbias pcasc net10[34] enb_10000_1 avss src_10000_1 bias_pstack
x10[33] avdd pbias pcasc net10[33] enb_10000_1 avss src_10000_1 bias_pstack
x10[32] avdd pbias pcasc net10[32] enb_10000_1 avss src_10000_1 bias_pstack
x10[31] avdd pbias pcasc net10[31] enb_10000_1 avss src_10000_1 bias_pstack
x10[30] avdd pbias pcasc net10[30] enb_10000_1 avss src_10000_1 bias_pstack
x10[29] avdd pbias pcasc net10[29] enb_10000_1 avss src_10000_1 bias_pstack
x10[28] avdd pbias pcasc net10[28] enb_10000_1 avss src_10000_1 bias_pstack
x10[27] avdd pbias pcasc net10[27] enb_10000_1 avss src_10000_1 bias_pstack
x10[26] avdd pbias pcasc net10[26] enb_10000_1 avss src_10000_1 bias_pstack
x10[25] avdd pbias pcasc net10[25] enb_10000_1 avss src_10000_1 bias_pstack
x10[24] avdd pbias pcasc net10[24] enb_10000_1 avss src_10000_1 bias_pstack
x10[23] avdd pbias pcasc net10[23] enb_10000_1 avss src_10000_1 bias_pstack
x10[22] avdd pbias pcasc net10[22] enb_10000_1 avss src_10000_1 bias_pstack
x10[21] avdd pbias pcasc net10[21] enb_10000_1 avss src_10000_1 bias_pstack
x10[20] avdd pbias pcasc net10[20] enb_10000_1 avss src_10000_1 bias_pstack
x10[19] avdd pbias pcasc net10[19] enb_10000_1 avss src_10000_1 bias_pstack
x10[18] avdd pbias pcasc net10[18] enb_10000_1 avss src_10000_1 bias_pstack
x10[17] avdd pbias pcasc net10[17] enb_10000_1 avss src_10000_1 bias_pstack
x10[16] avdd pbias pcasc net10[16] enb_10000_1 avss src_10000_1 bias_pstack
x10[15] avdd pbias pcasc net10[15] enb_10000_1 avss src_10000_1 bias_pstack
x10[14] avdd pbias pcasc net10[14] enb_10000_1 avss src_10000_1 bias_pstack
x10[13] avdd pbias pcasc net10[13] enb_10000_1 avss src_10000_1 bias_pstack
x10[12] avdd pbias pcasc net10[12] enb_10000_1 avss src_10000_1 bias_pstack
x10[11] avdd pbias pcasc net10[11] enb_10000_1 avss src_10000_1 bias_pstack
x10[10] avdd pbias pcasc net10[10] enb_10000_1 avss src_10000_1 bias_pstack
x10[9] avdd pbias pcasc net10[9] enb_10000_1 avss src_10000_1 bias_pstack
x10[8] avdd pbias pcasc net10[8] enb_10000_1 avss src_10000_1 bias_pstack
x10[7] avdd pbias pcasc net10[7] enb_10000_1 avss src_10000_1 bias_pstack
x10[6] avdd pbias pcasc net10[6] enb_10000_1 avss src_10000_1 bias_pstack
x10[5] avdd pbias pcasc net10[5] enb_10000_1 avss src_10000_1 bias_pstack
x10[4] avdd pbias pcasc net10[4] enb_10000_1 avss src_10000_1 bias_pstack
x10[3] avdd pbias pcasc net10[3] enb_10000_1 avss src_10000_1 bias_pstack
x10[2] avdd pbias pcasc net10[2] enb_10000_1 avss src_10000_1 bias_pstack
x10[1] avdd pbias pcasc net10[1] enb_10000_1 avss src_10000_1 bias_pstack
x10[0] avdd pbias pcasc net10[0] enb_10000_1 avss src_10000_1 bias_pstack
x1[99] snk_5000_1 ena_5000_1 net11[99] nbias avss bias_nstack
x1[98] snk_5000_1 ena_5000_1 net11[98] nbias avss bias_nstack
x1[97] snk_5000_1 ena_5000_1 net11[97] nbias avss bias_nstack
x1[96] snk_5000_1 ena_5000_1 net11[96] nbias avss bias_nstack
x1[95] snk_5000_1 ena_5000_1 net11[95] nbias avss bias_nstack
x1[94] snk_5000_1 ena_5000_1 net11[94] nbias avss bias_nstack
x1[93] snk_5000_1 ena_5000_1 net11[93] nbias avss bias_nstack
x1[92] snk_5000_1 ena_5000_1 net11[92] nbias avss bias_nstack
x1[91] snk_5000_1 ena_5000_1 net11[91] nbias avss bias_nstack
x1[90] snk_5000_1 ena_5000_1 net11[90] nbias avss bias_nstack
x1[89] snk_5000_1 ena_5000_1 net11[89] nbias avss bias_nstack
x1[88] snk_5000_1 ena_5000_1 net11[88] nbias avss bias_nstack
x1[87] snk_5000_1 ena_5000_1 net11[87] nbias avss bias_nstack
x1[86] snk_5000_1 ena_5000_1 net11[86] nbias avss bias_nstack
x1[85] snk_5000_1 ena_5000_1 net11[85] nbias avss bias_nstack
x1[84] snk_5000_1 ena_5000_1 net11[84] nbias avss bias_nstack
x1[83] snk_5000_1 ena_5000_1 net11[83] nbias avss bias_nstack
x1[82] snk_5000_1 ena_5000_1 net11[82] nbias avss bias_nstack
x1[81] snk_5000_1 ena_5000_1 net11[81] nbias avss bias_nstack
x1[80] snk_5000_1 ena_5000_1 net11[80] nbias avss bias_nstack
x1[79] snk_5000_1 ena_5000_1 net11[79] nbias avss bias_nstack
x1[78] snk_5000_1 ena_5000_1 net11[78] nbias avss bias_nstack
x1[77] snk_5000_1 ena_5000_1 net11[77] nbias avss bias_nstack
x1[76] snk_5000_1 ena_5000_1 net11[76] nbias avss bias_nstack
x1[75] snk_5000_1 ena_5000_1 net11[75] nbias avss bias_nstack
x1[74] snk_5000_1 ena_5000_1 net11[74] nbias avss bias_nstack
x1[73] snk_5000_1 ena_5000_1 net11[73] nbias avss bias_nstack
x1[72] snk_5000_1 ena_5000_1 net11[72] nbias avss bias_nstack
x1[71] snk_5000_1 ena_5000_1 net11[71] nbias avss bias_nstack
x1[70] snk_5000_1 ena_5000_1 net11[70] nbias avss bias_nstack
x1[69] snk_5000_1 ena_5000_1 net11[69] nbias avss bias_nstack
x1[68] snk_5000_1 ena_5000_1 net11[68] nbias avss bias_nstack
x1[67] snk_5000_1 ena_5000_1 net11[67] nbias avss bias_nstack
x1[66] snk_5000_1 ena_5000_1 net11[66] nbias avss bias_nstack
x1[65] snk_5000_1 ena_5000_1 net11[65] nbias avss bias_nstack
x1[64] snk_5000_1 ena_5000_1 net11[64] nbias avss bias_nstack
x1[63] snk_5000_1 ena_5000_1 net11[63] nbias avss bias_nstack
x1[62] snk_5000_1 ena_5000_1 net11[62] nbias avss bias_nstack
x1[61] snk_5000_1 ena_5000_1 net11[61] nbias avss bias_nstack
x1[60] snk_5000_1 ena_5000_1 net11[60] nbias avss bias_nstack
x1[59] snk_5000_1 ena_5000_1 net11[59] nbias avss bias_nstack
x1[58] snk_5000_1 ena_5000_1 net11[58] nbias avss bias_nstack
x1[57] snk_5000_1 ena_5000_1 net11[57] nbias avss bias_nstack
x1[56] snk_5000_1 ena_5000_1 net11[56] nbias avss bias_nstack
x1[55] snk_5000_1 ena_5000_1 net11[55] nbias avss bias_nstack
x1[54] snk_5000_1 ena_5000_1 net11[54] nbias avss bias_nstack
x1[53] snk_5000_1 ena_5000_1 net11[53] nbias avss bias_nstack
x1[52] snk_5000_1 ena_5000_1 net11[52] nbias avss bias_nstack
x1[51] snk_5000_1 ena_5000_1 net11[51] nbias avss bias_nstack
x1[50] snk_5000_1 ena_5000_1 net11[50] nbias avss bias_nstack
x1[49] snk_5000_1 ena_5000_1 net11[49] nbias avss bias_nstack
x1[48] snk_5000_1 ena_5000_1 net11[48] nbias avss bias_nstack
x1[47] snk_5000_1 ena_5000_1 net11[47] nbias avss bias_nstack
x1[46] snk_5000_1 ena_5000_1 net11[46] nbias avss bias_nstack
x1[45] snk_5000_1 ena_5000_1 net11[45] nbias avss bias_nstack
x1[44] snk_5000_1 ena_5000_1 net11[44] nbias avss bias_nstack
x1[43] snk_5000_1 ena_5000_1 net11[43] nbias avss bias_nstack
x1[42] snk_5000_1 ena_5000_1 net11[42] nbias avss bias_nstack
x1[41] snk_5000_1 ena_5000_1 net11[41] nbias avss bias_nstack
x1[40] snk_5000_1 ena_5000_1 net11[40] nbias avss bias_nstack
x1[39] snk_5000_1 ena_5000_1 net11[39] nbias avss bias_nstack
x1[38] snk_5000_1 ena_5000_1 net11[38] nbias avss bias_nstack
x1[37] snk_5000_1 ena_5000_1 net11[37] nbias avss bias_nstack
x1[36] snk_5000_1 ena_5000_1 net11[36] nbias avss bias_nstack
x1[35] snk_5000_1 ena_5000_1 net11[35] nbias avss bias_nstack
x1[34] snk_5000_1 ena_5000_1 net11[34] nbias avss bias_nstack
x1[33] snk_5000_1 ena_5000_1 net11[33] nbias avss bias_nstack
x1[32] snk_5000_1 ena_5000_1 net11[32] nbias avss bias_nstack
x1[31] snk_5000_1 ena_5000_1 net11[31] nbias avss bias_nstack
x1[30] snk_5000_1 ena_5000_1 net11[30] nbias avss bias_nstack
x1[29] snk_5000_1 ena_5000_1 net11[29] nbias avss bias_nstack
x1[28] snk_5000_1 ena_5000_1 net11[28] nbias avss bias_nstack
x1[27] snk_5000_1 ena_5000_1 net11[27] nbias avss bias_nstack
x1[26] snk_5000_1 ena_5000_1 net11[26] nbias avss bias_nstack
x1[25] snk_5000_1 ena_5000_1 net11[25] nbias avss bias_nstack
x1[24] snk_5000_1 ena_5000_1 net11[24] nbias avss bias_nstack
x1[23] snk_5000_1 ena_5000_1 net11[23] nbias avss bias_nstack
x1[22] snk_5000_1 ena_5000_1 net11[22] nbias avss bias_nstack
x1[21] snk_5000_1 ena_5000_1 net11[21] nbias avss bias_nstack
x1[20] snk_5000_1 ena_5000_1 net11[20] nbias avss bias_nstack
x1[19] snk_5000_1 ena_5000_1 net11[19] nbias avss bias_nstack
x1[18] snk_5000_1 ena_5000_1 net11[18] nbias avss bias_nstack
x1[17] snk_5000_1 ena_5000_1 net11[17] nbias avss bias_nstack
x1[16] snk_5000_1 ena_5000_1 net11[16] nbias avss bias_nstack
x1[15] snk_5000_1 ena_5000_1 net11[15] nbias avss bias_nstack
x1[14] snk_5000_1 ena_5000_1 net11[14] nbias avss bias_nstack
x1[13] snk_5000_1 ena_5000_1 net11[13] nbias avss bias_nstack
x1[12] snk_5000_1 ena_5000_1 net11[12] nbias avss bias_nstack
x1[11] snk_5000_1 ena_5000_1 net11[11] nbias avss bias_nstack
x1[10] snk_5000_1 ena_5000_1 net11[10] nbias avss bias_nstack
x1[9] snk_5000_1 ena_5000_1 net11[9] nbias avss bias_nstack
x1[8] snk_5000_1 ena_5000_1 net11[8] nbias avss bias_nstack
x1[7] snk_5000_1 ena_5000_1 net11[7] nbias avss bias_nstack
x1[6] snk_5000_1 ena_5000_1 net11[6] nbias avss bias_nstack
x1[5] snk_5000_1 ena_5000_1 net11[5] nbias avss bias_nstack
x1[4] snk_5000_1 ena_5000_1 net11[4] nbias avss bias_nstack
x1[3] snk_5000_1 ena_5000_1 net11[3] nbias avss bias_nstack
x1[2] snk_5000_1 ena_5000_1 net11[2] nbias avss bias_nstack
x1[1] snk_5000_1 ena_5000_1 net11[1] nbias avss bias_nstack
x1[0] snk_5000_1 ena_5000_1 net11[0] nbias avss bias_nstack
x3[99] snk_5000_2 ena_5000_2 net12[99] nbias avss bias_nstack
x3[98] snk_5000_2 ena_5000_2 net12[98] nbias avss bias_nstack
x3[97] snk_5000_2 ena_5000_2 net12[97] nbias avss bias_nstack
x3[96] snk_5000_2 ena_5000_2 net12[96] nbias avss bias_nstack
x3[95] snk_5000_2 ena_5000_2 net12[95] nbias avss bias_nstack
x3[94] snk_5000_2 ena_5000_2 net12[94] nbias avss bias_nstack
x3[93] snk_5000_2 ena_5000_2 net12[93] nbias avss bias_nstack
x3[92] snk_5000_2 ena_5000_2 net12[92] nbias avss bias_nstack
x3[91] snk_5000_2 ena_5000_2 net12[91] nbias avss bias_nstack
x3[90] snk_5000_2 ena_5000_2 net12[90] nbias avss bias_nstack
x3[89] snk_5000_2 ena_5000_2 net12[89] nbias avss bias_nstack
x3[88] snk_5000_2 ena_5000_2 net12[88] nbias avss bias_nstack
x3[87] snk_5000_2 ena_5000_2 net12[87] nbias avss bias_nstack
x3[86] snk_5000_2 ena_5000_2 net12[86] nbias avss bias_nstack
x3[85] snk_5000_2 ena_5000_2 net12[85] nbias avss bias_nstack
x3[84] snk_5000_2 ena_5000_2 net12[84] nbias avss bias_nstack
x3[83] snk_5000_2 ena_5000_2 net12[83] nbias avss bias_nstack
x3[82] snk_5000_2 ena_5000_2 net12[82] nbias avss bias_nstack
x3[81] snk_5000_2 ena_5000_2 net12[81] nbias avss bias_nstack
x3[80] snk_5000_2 ena_5000_2 net12[80] nbias avss bias_nstack
x3[79] snk_5000_2 ena_5000_2 net12[79] nbias avss bias_nstack
x3[78] snk_5000_2 ena_5000_2 net12[78] nbias avss bias_nstack
x3[77] snk_5000_2 ena_5000_2 net12[77] nbias avss bias_nstack
x3[76] snk_5000_2 ena_5000_2 net12[76] nbias avss bias_nstack
x3[75] snk_5000_2 ena_5000_2 net12[75] nbias avss bias_nstack
x3[74] snk_5000_2 ena_5000_2 net12[74] nbias avss bias_nstack
x3[73] snk_5000_2 ena_5000_2 net12[73] nbias avss bias_nstack
x3[72] snk_5000_2 ena_5000_2 net12[72] nbias avss bias_nstack
x3[71] snk_5000_2 ena_5000_2 net12[71] nbias avss bias_nstack
x3[70] snk_5000_2 ena_5000_2 net12[70] nbias avss bias_nstack
x3[69] snk_5000_2 ena_5000_2 net12[69] nbias avss bias_nstack
x3[68] snk_5000_2 ena_5000_2 net12[68] nbias avss bias_nstack
x3[67] snk_5000_2 ena_5000_2 net12[67] nbias avss bias_nstack
x3[66] snk_5000_2 ena_5000_2 net12[66] nbias avss bias_nstack
x3[65] snk_5000_2 ena_5000_2 net12[65] nbias avss bias_nstack
x3[64] snk_5000_2 ena_5000_2 net12[64] nbias avss bias_nstack
x3[63] snk_5000_2 ena_5000_2 net12[63] nbias avss bias_nstack
x3[62] snk_5000_2 ena_5000_2 net12[62] nbias avss bias_nstack
x3[61] snk_5000_2 ena_5000_2 net12[61] nbias avss bias_nstack
x3[60] snk_5000_2 ena_5000_2 net12[60] nbias avss bias_nstack
x3[59] snk_5000_2 ena_5000_2 net12[59] nbias avss bias_nstack
x3[58] snk_5000_2 ena_5000_2 net12[58] nbias avss bias_nstack
x3[57] snk_5000_2 ena_5000_2 net12[57] nbias avss bias_nstack
x3[56] snk_5000_2 ena_5000_2 net12[56] nbias avss bias_nstack
x3[55] snk_5000_2 ena_5000_2 net12[55] nbias avss bias_nstack
x3[54] snk_5000_2 ena_5000_2 net12[54] nbias avss bias_nstack
x3[53] snk_5000_2 ena_5000_2 net12[53] nbias avss bias_nstack
x3[52] snk_5000_2 ena_5000_2 net12[52] nbias avss bias_nstack
x3[51] snk_5000_2 ena_5000_2 net12[51] nbias avss bias_nstack
x3[50] snk_5000_2 ena_5000_2 net12[50] nbias avss bias_nstack
x3[49] snk_5000_2 ena_5000_2 net12[49] nbias avss bias_nstack
x3[48] snk_5000_2 ena_5000_2 net12[48] nbias avss bias_nstack
x3[47] snk_5000_2 ena_5000_2 net12[47] nbias avss bias_nstack
x3[46] snk_5000_2 ena_5000_2 net12[46] nbias avss bias_nstack
x3[45] snk_5000_2 ena_5000_2 net12[45] nbias avss bias_nstack
x3[44] snk_5000_2 ena_5000_2 net12[44] nbias avss bias_nstack
x3[43] snk_5000_2 ena_5000_2 net12[43] nbias avss bias_nstack
x3[42] snk_5000_2 ena_5000_2 net12[42] nbias avss bias_nstack
x3[41] snk_5000_2 ena_5000_2 net12[41] nbias avss bias_nstack
x3[40] snk_5000_2 ena_5000_2 net12[40] nbias avss bias_nstack
x3[39] snk_5000_2 ena_5000_2 net12[39] nbias avss bias_nstack
x3[38] snk_5000_2 ena_5000_2 net12[38] nbias avss bias_nstack
x3[37] snk_5000_2 ena_5000_2 net12[37] nbias avss bias_nstack
x3[36] snk_5000_2 ena_5000_2 net12[36] nbias avss bias_nstack
x3[35] snk_5000_2 ena_5000_2 net12[35] nbias avss bias_nstack
x3[34] snk_5000_2 ena_5000_2 net12[34] nbias avss bias_nstack
x3[33] snk_5000_2 ena_5000_2 net12[33] nbias avss bias_nstack
x3[32] snk_5000_2 ena_5000_2 net12[32] nbias avss bias_nstack
x3[31] snk_5000_2 ena_5000_2 net12[31] nbias avss bias_nstack
x3[30] snk_5000_2 ena_5000_2 net12[30] nbias avss bias_nstack
x3[29] snk_5000_2 ena_5000_2 net12[29] nbias avss bias_nstack
x3[28] snk_5000_2 ena_5000_2 net12[28] nbias avss bias_nstack
x3[27] snk_5000_2 ena_5000_2 net12[27] nbias avss bias_nstack
x3[26] snk_5000_2 ena_5000_2 net12[26] nbias avss bias_nstack
x3[25] snk_5000_2 ena_5000_2 net12[25] nbias avss bias_nstack
x3[24] snk_5000_2 ena_5000_2 net12[24] nbias avss bias_nstack
x3[23] snk_5000_2 ena_5000_2 net12[23] nbias avss bias_nstack
x3[22] snk_5000_2 ena_5000_2 net12[22] nbias avss bias_nstack
x3[21] snk_5000_2 ena_5000_2 net12[21] nbias avss bias_nstack
x3[20] snk_5000_2 ena_5000_2 net12[20] nbias avss bias_nstack
x3[19] snk_5000_2 ena_5000_2 net12[19] nbias avss bias_nstack
x3[18] snk_5000_2 ena_5000_2 net12[18] nbias avss bias_nstack
x3[17] snk_5000_2 ena_5000_2 net12[17] nbias avss bias_nstack
x3[16] snk_5000_2 ena_5000_2 net12[16] nbias avss bias_nstack
x3[15] snk_5000_2 ena_5000_2 net12[15] nbias avss bias_nstack
x3[14] snk_5000_2 ena_5000_2 net12[14] nbias avss bias_nstack
x3[13] snk_5000_2 ena_5000_2 net12[13] nbias avss bias_nstack
x3[12] snk_5000_2 ena_5000_2 net12[12] nbias avss bias_nstack
x3[11] snk_5000_2 ena_5000_2 net12[11] nbias avss bias_nstack
x3[10] snk_5000_2 ena_5000_2 net12[10] nbias avss bias_nstack
x3[9] snk_5000_2 ena_5000_2 net12[9] nbias avss bias_nstack
x3[8] snk_5000_2 ena_5000_2 net12[8] nbias avss bias_nstack
x3[7] snk_5000_2 ena_5000_2 net12[7] nbias avss bias_nstack
x3[6] snk_5000_2 ena_5000_2 net12[6] nbias avss bias_nstack
x3[5] snk_5000_2 ena_5000_2 net12[5] nbias avss bias_nstack
x3[4] snk_5000_2 ena_5000_2 net12[4] nbias avss bias_nstack
x3[3] snk_5000_2 ena_5000_2 net12[3] nbias avss bias_nstack
x3[2] snk_5000_2 ena_5000_2 net12[2] nbias avss bias_nstack
x3[1] snk_5000_2 ena_5000_2 net12[1] nbias avss bias_nstack
x3[0] snk_5000_2 ena_5000_2 net12[0] nbias avss bias_nstack
x4[11] avdd pbias pcasc net13[11] enb_600 avss src_600 bias_pstack
x4[10] avdd pbias pcasc net13[10] enb_600 avss src_600 bias_pstack
x4[9] avdd pbias pcasc net13[9] enb_600 avss src_600 bias_pstack
x4[8] avdd pbias pcasc net13[8] enb_600 avss src_600 bias_pstack
x4[7] avdd pbias pcasc net13[7] enb_600 avss src_600 bias_pstack
x4[6] avdd pbias pcasc net13[6] enb_600 avss src_600 bias_pstack
x4[5] avdd pbias pcasc net13[5] enb_600 avss src_600 bias_pstack
x4[4] avdd pbias pcasc net13[4] enb_600 avss src_600 bias_pstack
x4[3] avdd pbias pcasc net13[3] enb_600 avss src_600 bias_pstack
x4[2] avdd pbias pcasc net13[2] enb_600 avss src_600 bias_pstack
x4[1] avdd pbias pcasc net13[1] enb_600 avss src_600 bias_pstack
x4[0] avdd pbias pcasc net13[0] enb_600 avss src_600 bias_pstack
x5[7] avdd pbias pcasc net14[7] enb_400 avss src_400 bias_pstack
x5[6] avdd pbias pcasc net14[6] enb_400 avss src_400 bias_pstack
x5[5] avdd pbias pcasc net14[5] enb_400 avss src_400 bias_pstack
x5[4] avdd pbias pcasc net14[4] enb_400 avss src_400 bias_pstack
x5[3] avdd pbias pcasc net14[3] enb_400 avss src_400 bias_pstack
x5[2] avdd pbias pcasc net14[2] enb_400 avss src_400 bias_pstack
x5[1] avdd pbias pcasc net14[1] enb_400 avss src_400 bias_pstack
x5[0] avdd pbias pcasc net14[0] enb_400 avss src_400 bias_pstack
x6[3] avdd pbias pcasc net15[3] enb_200_0 avss src_200_0 bias_pstack
x6[2] avdd pbias pcasc net15[2] enb_200_0 avss src_200_0 bias_pstack
x6[1] avdd pbias pcasc net15[1] enb_200_0 avss src_200_0 bias_pstack
x6[0] avdd pbias pcasc net15[0] enb_200_0 avss src_200_0 bias_pstack
x7[3] avdd pbias pcasc net16[3] enb_200_1 avss src_200_1 bias_pstack
x7[2] avdd pbias pcasc net16[2] enb_200_1 avss src_200_1 bias_pstack
x7[1] avdd pbias pcasc net16[1] enb_200_1 avss src_200_1 bias_pstack
x7[0] avdd pbias pcasc net16[0] enb_200_1 avss src_200_1 bias_pstack
x11[3] avdd pbias pcasc net17[3] enb_200_2 avss src_200_2 bias_pstack
x11[2] avdd pbias pcasc net17[2] enb_200_2 avss src_200_2 bias_pstack
x11[1] avdd pbias pcasc net17[1] enb_200_2 avss src_200_2 bias_pstack
x11[0] avdd pbias pcasc net17[0] enb_200_2 avss src_200_2 bias_pstack
x12[1] avdd pbias pcasc net18[1] enb_100 avss src_100 bias_pstack
x12[0] avdd pbias pcasc net18[0] enb_100 avss src_100 bias_pstack
x13 avdd pbias pcasc net19 enb_50 avss src_50 bias_pstack
x14[74] snk_3700 ena_3700 net20[74] nbias avss bias_nstack
x14[73] snk_3700 ena_3700 net20[73] nbias avss bias_nstack
x14[72] snk_3700 ena_3700 net20[72] nbias avss bias_nstack
x14[71] snk_3700 ena_3700 net20[71] nbias avss bias_nstack
x14[70] snk_3700 ena_3700 net20[70] nbias avss bias_nstack
x14[69] snk_3700 ena_3700 net20[69] nbias avss bias_nstack
x14[68] snk_3700 ena_3700 net20[68] nbias avss bias_nstack
x14[67] snk_3700 ena_3700 net20[67] nbias avss bias_nstack
x14[66] snk_3700 ena_3700 net20[66] nbias avss bias_nstack
x14[65] snk_3700 ena_3700 net20[65] nbias avss bias_nstack
x14[64] snk_3700 ena_3700 net20[64] nbias avss bias_nstack
x14[63] snk_3700 ena_3700 net20[63] nbias avss bias_nstack
x14[62] snk_3700 ena_3700 net20[62] nbias avss bias_nstack
x14[61] snk_3700 ena_3700 net20[61] nbias avss bias_nstack
x14[60] snk_3700 ena_3700 net20[60] nbias avss bias_nstack
x14[59] snk_3700 ena_3700 net20[59] nbias avss bias_nstack
x14[58] snk_3700 ena_3700 net20[58] nbias avss bias_nstack
x14[57] snk_3700 ena_3700 net20[57] nbias avss bias_nstack
x14[56] snk_3700 ena_3700 net20[56] nbias avss bias_nstack
x14[55] snk_3700 ena_3700 net20[55] nbias avss bias_nstack
x14[54] snk_3700 ena_3700 net20[54] nbias avss bias_nstack
x14[53] snk_3700 ena_3700 net20[53] nbias avss bias_nstack
x14[52] snk_3700 ena_3700 net20[52] nbias avss bias_nstack
x14[51] snk_3700 ena_3700 net20[51] nbias avss bias_nstack
x14[50] snk_3700 ena_3700 net20[50] nbias avss bias_nstack
x14[49] snk_3700 ena_3700 net20[49] nbias avss bias_nstack
x14[48] snk_3700 ena_3700 net20[48] nbias avss bias_nstack
x14[47] snk_3700 ena_3700 net20[47] nbias avss bias_nstack
x14[46] snk_3700 ena_3700 net20[46] nbias avss bias_nstack
x14[45] snk_3700 ena_3700 net20[45] nbias avss bias_nstack
x14[44] snk_3700 ena_3700 net20[44] nbias avss bias_nstack
x14[43] snk_3700 ena_3700 net20[43] nbias avss bias_nstack
x14[42] snk_3700 ena_3700 net20[42] nbias avss bias_nstack
x14[41] snk_3700 ena_3700 net20[41] nbias avss bias_nstack
x14[40] snk_3700 ena_3700 net20[40] nbias avss bias_nstack
x14[39] snk_3700 ena_3700 net20[39] nbias avss bias_nstack
x14[38] snk_3700 ena_3700 net20[38] nbias avss bias_nstack
x14[37] snk_3700 ena_3700 net20[37] nbias avss bias_nstack
x14[36] snk_3700 ena_3700 net20[36] nbias avss bias_nstack
x14[35] snk_3700 ena_3700 net20[35] nbias avss bias_nstack
x14[34] snk_3700 ena_3700 net20[34] nbias avss bias_nstack
x14[33] snk_3700 ena_3700 net20[33] nbias avss bias_nstack
x14[32] snk_3700 ena_3700 net20[32] nbias avss bias_nstack
x14[31] snk_3700 ena_3700 net20[31] nbias avss bias_nstack
x14[30] snk_3700 ena_3700 net20[30] nbias avss bias_nstack
x14[29] snk_3700 ena_3700 net20[29] nbias avss bias_nstack
x14[28] snk_3700 ena_3700 net20[28] nbias avss bias_nstack
x14[27] snk_3700 ena_3700 net20[27] nbias avss bias_nstack
x14[26] snk_3700 ena_3700 net20[26] nbias avss bias_nstack
x14[25] snk_3700 ena_3700 net20[25] nbias avss bias_nstack
x14[24] snk_3700 ena_3700 net20[24] nbias avss bias_nstack
x14[23] snk_3700 ena_3700 net20[23] nbias avss bias_nstack
x14[22] snk_3700 ena_3700 net20[22] nbias avss bias_nstack
x14[21] snk_3700 ena_3700 net20[21] nbias avss bias_nstack
x14[20] snk_3700 ena_3700 net20[20] nbias avss bias_nstack
x14[19] snk_3700 ena_3700 net20[19] nbias avss bias_nstack
x14[18] snk_3700 ena_3700 net20[18] nbias avss bias_nstack
x14[17] snk_3700 ena_3700 net20[17] nbias avss bias_nstack
x14[16] snk_3700 ena_3700 net20[16] nbias avss bias_nstack
x14[15] snk_3700 ena_3700 net20[15] nbias avss bias_nstack
x14[14] snk_3700 ena_3700 net20[14] nbias avss bias_nstack
x14[13] snk_3700 ena_3700 net20[13] nbias avss bias_nstack
x14[12] snk_3700 ena_3700 net20[12] nbias avss bias_nstack
x14[11] snk_3700 ena_3700 net20[11] nbias avss bias_nstack
x14[10] snk_3700 ena_3700 net20[10] nbias avss bias_nstack
x14[9] snk_3700 ena_3700 net20[9] nbias avss bias_nstack
x14[8] snk_3700 ena_3700 net20[8] nbias avss bias_nstack
x14[7] snk_3700 ena_3700 net20[7] nbias avss bias_nstack
x14[6] snk_3700 ena_3700 net20[6] nbias avss bias_nstack
x14[5] snk_3700 ena_3700 net20[5] nbias avss bias_nstack
x14[4] snk_3700 ena_3700 net20[4] nbias avss bias_nstack
x14[3] snk_3700 ena_3700 net20[3] nbias avss bias_nstack
x14[2] snk_3700 ena_3700 net20[2] nbias avss bias_nstack
x14[1] snk_3700 ena_3700 net20[1] nbias avss bias_nstack
x14[0] snk_3700 ena_3700 net20[0] nbias avss bias_nstack
x15[39] snk_2000 ena_2000 net21[39] nbias avss bias_nstack
x15[38] snk_2000 ena_2000 net21[38] nbias avss bias_nstack
x15[37] snk_2000 ena_2000 net21[37] nbias avss bias_nstack
x15[36] snk_2000 ena_2000 net21[36] nbias avss bias_nstack
x15[35] snk_2000 ena_2000 net21[35] nbias avss bias_nstack
x15[34] snk_2000 ena_2000 net21[34] nbias avss bias_nstack
x15[33] snk_2000 ena_2000 net21[33] nbias avss bias_nstack
x15[32] snk_2000 ena_2000 net21[32] nbias avss bias_nstack
x15[31] snk_2000 ena_2000 net21[31] nbias avss bias_nstack
x15[30] snk_2000 ena_2000 net21[30] nbias avss bias_nstack
x15[29] snk_2000 ena_2000 net21[29] nbias avss bias_nstack
x15[28] snk_2000 ena_2000 net21[28] nbias avss bias_nstack
x15[27] snk_2000 ena_2000 net21[27] nbias avss bias_nstack
x15[26] snk_2000 ena_2000 net21[26] nbias avss bias_nstack
x15[25] snk_2000 ena_2000 net21[25] nbias avss bias_nstack
x15[24] snk_2000 ena_2000 net21[24] nbias avss bias_nstack
x15[23] snk_2000 ena_2000 net21[23] nbias avss bias_nstack
x15[22] snk_2000 ena_2000 net21[22] nbias avss bias_nstack
x15[21] snk_2000 ena_2000 net21[21] nbias avss bias_nstack
x15[20] snk_2000 ena_2000 net21[20] nbias avss bias_nstack
x15[19] snk_2000 ena_2000 net21[19] nbias avss bias_nstack
x15[18] snk_2000 ena_2000 net21[18] nbias avss bias_nstack
x15[17] snk_2000 ena_2000 net21[17] nbias avss bias_nstack
x15[16] snk_2000 ena_2000 net21[16] nbias avss bias_nstack
x15[15] snk_2000 ena_2000 net21[15] nbias avss bias_nstack
x15[14] snk_2000 ena_2000 net21[14] nbias avss bias_nstack
x15[13] snk_2000 ena_2000 net21[13] nbias avss bias_nstack
x15[12] snk_2000 ena_2000 net21[12] nbias avss bias_nstack
x15[11] snk_2000 ena_2000 net21[11] nbias avss bias_nstack
x15[10] snk_2000 ena_2000 net21[10] nbias avss bias_nstack
x15[9] snk_2000 ena_2000 net21[9] nbias avss bias_nstack
x15[8] snk_2000 ena_2000 net21[8] nbias avss bias_nstack
x15[7] snk_2000 ena_2000 net21[7] nbias avss bias_nstack
x15[6] snk_2000 ena_2000 net21[6] nbias avss bias_nstack
x15[5] snk_2000 ena_2000 net21[5] nbias avss bias_nstack
x15[4] snk_2000 ena_2000 net21[4] nbias avss bias_nstack
x15[3] snk_2000 ena_2000 net21[3] nbias avss bias_nstack
x15[2] snk_2000 ena_2000 net21[2] nbias avss bias_nstack
x15[1] snk_2000 ena_2000 net21[1] nbias avss bias_nstack
x15[0] snk_2000 ena_2000 net21[0] nbias avss bias_nstack
.ends


* expanding   symbol:  power_stage.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/power_stage.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/power_stage.sch
.subckt power_stage P_IN P_IN_N VSS VDD_PWR SW_NODE
*.PININFO P_IN:I P_IN_N:I SW_NODE:I VDD_PWR:I VSS:I
XM14 SW_NODE P_DRIVE VDD_PWR VDD_PWR sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4.38 nf=1 m=4512
x2 P_IN P_IN_N VDD_PWR VSS P_DRIVE gate_drive
.ends


* expanding   symbol:  chipalooza/lpopamp.sym # of pins=9
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/lpopamp.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/lpopamp.sch
.subckt lpopamp im o ib vsub avss avdd enb en ip

.ends


* expanding   symbol:  chipalooza/sky130_ajc_ip__brownout.sym # of pins=22
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ajc_ip__brownout.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ajc_ip__brownout.sch
.subckt sky130_ajc_ip__brownout avdd avss outb dvdd osc_ck dvss dcomp vbg_1v2 otrip[2] otrip[1] otrip[0] itest brout_filt vtrip[2]
+ vtrip[1] vtrip[0] vin_brout ena force_ena_rc_osc vin_vunder force_dis_rc_osc timed_out vunder force_short_oneshot isrc_sel ibg_200n

.ends


* expanding   symbol:  chipalooza/sky130_ajc_ip__overvoltage.sym # of pins=12
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ajc_ip__overvoltage.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ajc_ip__overvoltage.sch
.subckt sky130_ajc_ip__overvoltage avdd avss dvdd dvss vbg_1v2 ovout itest otrip[3] otrip[2] otrip[1] otrip[0] vin ena isrc_sel
+ ibg_200n

.ends


* expanding   symbol:  chipalooza/sky130_ajc_ip__por.sym # of pins=22
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ajc_ip__por.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ajc_ip__por.sch
.subckt sky130_ajc_ip__por avdd porb_h porb avss dvdd por dvss osc_ck vbg_1v2 dcomp otrip[2] otrip[1] otrip[0] itest force_pdn
+ pwup_filt vin force_ena_rc_osc force_dis_rc_osc startup_timed_out por_timed_out force_short_oneshot isrc_sel ibg_200n

.ends


* expanding   symbol:  chipalooza/sky130_ak_ip__comparator.sym # of pins=10
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ak_ip__comparator.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ak_ip__comparator.sch
.subckt sky130_ak_ip__comparator DVDD AVDD AGND Vinp Vout Vinm en hyst[1] hyst[0] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0]
+ ibias

.ends


* expanding   symbol:  chipalooza/sky130_be_ip__lsxo.sym # of pins=10
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_be_ip__lsxo.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_be_ip__lsxo.sch
.subckt sky130_be_ip__lsxo avdd avss dvdd dvss ibias ena standby dout xin xout

.ends


* expanding   symbol:  chipalooza/sky130_ht_ip__hsxo_cpz1.sym # of pins=11
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ht_ip__hsxo_cpz1.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_ht_ip__hsxo_cpz1.sch
.subckt sky130_ht_ip__hsxo_cpz1 XOUT XIN ENA STDBY DOUT AVDD DVDD AVSS DVSS IBIAS GUARD

.ends


* expanding   symbol:  chipalooza/sky130_td_ip__opamp_hp.sym # of pins=9
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_td_ip__opamp_hp.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_td_ip__opamp_hp.sch
.subckt sky130_td_ip__opamp_hp avdd vout ibias vinn vinp avss dvdd dvss ena

.ends


* expanding   symbol:  chipalooza/sky130_vbl_ip__overvoltage.sym # of pins=12
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_vbl_ip__overvoltage.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_vbl_ip__overvoltage.sch
.subckt sky130_vbl_ip__overvoltage avdd dvdd ena vtrip[3] ibias vtrip[2] ovout vbg vtrip[1] vtrip[0] dvss avss

.ends


* expanding   symbol:  lvl_shift_invert.sym # of pins=6
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/lvl_shift_invert.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/lvl_shift_invert.sch
.subckt lvl_shift_invert in1v8 out3v3 outb3v3 dvdd dvss avdd
*.PININFO in1v8:I dvdd:B dvss:B avdd:B out3v3:O outb3v3:O
x2 in1v8 dvdd dvss dvss avdd avdd out3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x4 out3v3 dvss dvss avdd avdd outb3v3 sky130_fd_sc_hvl__inv_2
.ends


* expanding   symbol:  analog_mux_sel1v8.sym # of pins=8
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/analog_mux_sel1v8.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/analog_mux_sel1v8.sch
.subckt analog_mux_sel1v8 avss selA inA avdd inB out dvdd dvss
*.PININFO selA:I avss:B out:B inA:B avdd:B inB:B dvdd:B dvss:B
x1 net1 avss inA out avdd isolated_switch
x2 selA dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
x3 net2 avss inB out avdd isolated_switch
x4 net1 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
.ends


* expanding   symbol:  isolated_switch_ena1v8.sym # of pins=7
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/isolated_switch_ena1v8.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/isolated_switch_ena1v8.sch
.subckt isolated_switch_ena1v8 dvdd dvss avss on out in avdd
*.PININFO on:I avss:B out:B in:B avdd:B
x1 net1 avss out in avdd isolated_switch
x2 on dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
.ends


* expanding   symbol:  chipalooza/sky130_od_ip__tempsensor_ext_vp.sym # of pins=6
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_od_ip__tempsensor_ext_vp.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/chipalooza/sky130_od_ip__tempsensor_ext_vp.sch
.subckt sky130_od_ip__tempsensor_ext_vp vbe1_out vdd vss vbg ena vbe2_out

.ends


* expanding   symbol:  weiser/bandgap.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/weiser/bandgap.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/weiser/bandgap.sch
.subckt bandgap vdd vbg vss bias trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7] trim[6] trim[5]
+ trim[4] trim[3] trim[2] trim[1] trim[0]

.ends


* expanding   symbol:  weiser/bias_basis_current.sym # of pins=4
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/weiser/bias_basis_current.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/weiser/bias_basis_current.sch
.subckt bias_basis_current vdd vss ibp ibn

.ends


* expanding   symbol:  bias_nstack.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/bias_nstack.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/bias_nstack.sch
.subckt bias_nstack itail ena vcasc nbias avss
*.PININFO avss:B ena:I nbias:I itail:B vcasc:B
XM3 net1 nbias avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XM6 vcasc nbias net1 avss sky130_fd_pr__nfet_05v0_nvt L=1 W=3 nf=1 m=1
XM12 itail ena vcasc avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XD1 avss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  bias_pstack.sym # of pins=7
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/bias_pstack.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/bias_pstack.sch
.subckt bias_pstack avdd pbias pcasc vcasc enb avss itail
*.PININFO avdd:B itail:B enb:I pcasc:I vcasc:B pbias:I avss:B
XM13 net1 pbias avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XM18 itail enb vcasc avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XM14 vcasc pcasc net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XD1 avss enb sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  gate_drive.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/gate_drive.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/gate_drive.sch
.subckt gate_drive IN_P IN_M VDD VSS OUT
*.PININFO IN_M:I IN_P:I VDD:I VSS:I OUT:O
XM1 net1 IN_P VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM2 net1 S1_N VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM3 S1_N IN_M VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM4 S1_N net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM5 S2_N S1_N VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 m=2
XM6 S2_N S1_N VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=2
XM7 S3_N S2_N VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 m=6
XM8 S3_N S2_N VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=6
XM9 S4_N S3_N VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 m=20
XM10 S4_N S3_N VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=20
XM11 OUT S4_N VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 m=60
XM12 OUT S4_N VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=60
.ends


* expanding   symbol:  isolated_switch.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_1/xschem/isolated_switch.sym
** sch_path: /home/tim/gits/chipalooza_projects_1/xschem/isolated_switch.sch
.subckt isolated_switch on vss out in vdd
*.PININFO on:I out:B vdd:B vss:B in:B
XM1 in onp net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=2 m=1
XM2 in onb net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM3 net1 onb net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM4 net1 onp net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM5 in onb in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM6 in onp in vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM7 onb on vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM8 onb on vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM9 onp onb vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM10 onp onb vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XXD1 vss on sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
XM11 net1 onp out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8 nf=2 m=1
XM12 net1 onb out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM13 out onb out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM14 out onp out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM15 net1 onb net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM16 net1 onp net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM17 vss onb net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends

.end
