magic
tech sky130A
magscale 1 2
timestamp 1714671808
<< locali >>
rect -21956 -11267 -14626 -11266
rect -22251 -11286 -14626 -11267
rect -22251 -11448 -14401 -11286
rect -22251 -29751 -22182 -11448
rect -22048 -11650 -14401 -11448
rect -22048 -12586 -21524 -11650
rect -16167 -12586 -14401 -11650
rect -22048 -12795 -14401 -12586
rect -22048 -12943 -14586 -12795
rect -22048 -29751 -21918 -12943
rect -22251 -29826 -21918 -29751
rect -14653 -29752 -14586 -12943
rect -14468 -29752 -14401 -12795
rect -14653 -29821 -14401 -29752
<< viali >>
rect -22182 -29751 -22048 -11448
rect -21524 -12586 -16167 -11650
rect -14586 -29752 -14468 -12795
rect -16687 -31085 -16653 -30895
rect -16603 -31007 -16281 -30973
rect -16137 -31083 -16103 -30893
rect -16050 -31007 -15733 -30973
rect -15679 -31006 -15558 -30971
<< metal1 >>
rect -14656 -11277 -11060 -11251
rect -21930 -11290 -11060 -11282
rect -22352 -11302 -11060 -11290
rect -86481 -11448 -11060 -11302
rect -86481 -12297 -22182 -11448
rect -85199 -28067 -79389 -13362
rect -78189 -28067 -67389 -13362
rect -66189 -28067 -55389 -13362
rect -54189 -28067 -43389 -13362
rect -42189 -28067 -31389 -13362
rect -30189 -28067 -23576 -13362
rect -85199 -30024 -23576 -28067
rect -22352 -29751 -22182 -12297
rect -22048 -11650 -11060 -11448
rect -22048 -12586 -21524 -11650
rect -16167 -12586 -11060 -11650
rect -22048 -12795 -11060 -12586
rect -22048 -12888 -14586 -12795
rect -22048 -29751 -21879 -12888
rect -21510 -29400 -21500 -13300
rect -21160 -29400 -21150 -13300
rect -15450 -29400 -15440 -13300
rect -15100 -29400 -15090 -13300
rect -85209 -32280 -85199 -30024
rect -23576 -32280 -23566 -30024
rect -22352 -31185 -21879 -29751
rect -14681 -29752 -14586 -12888
rect -14468 -12888 -11060 -12795
rect -14468 -29752 -13989 -12888
rect -14681 -29823 -13989 -29752
rect -17198 -30733 -11477 -30254
rect -16712 -30885 -16647 -30882
rect -16712 -31086 -16706 -30885
rect -16653 -31086 -16647 -30885
rect -16154 -30886 -16097 -30878
rect -16154 -30967 -16152 -30886
rect -16616 -30973 -16152 -30967
rect -16616 -31007 -16603 -30973
rect -16281 -31007 -16152 -30973
rect -16616 -31013 -16152 -31007
rect -16712 -31100 -16647 -31086
rect -16154 -31087 -16152 -31013
rect -16099 -31087 -16097 -30886
rect -16062 -30971 -15541 -30965
rect -16062 -30973 -15679 -30971
rect -16062 -31007 -16050 -30973
rect -15733 -31006 -15679 -30973
rect -15558 -31006 -15541 -30971
rect -15733 -31007 -15541 -31006
rect -16062 -31014 -15983 -31007
rect -15993 -31034 -15983 -31014
rect -15773 -31014 -15541 -31007
rect -15773 -31034 -15763 -31014
rect -15993 -31041 -15763 -31034
rect -16154 -31096 -16097 -31087
rect -22352 -31663 -15070 -31185
rect -22229 -31664 -15070 -31663
<< via1 >>
rect -21500 -29400 -21160 -13300
rect -15440 -29400 -15100 -13300
rect -85199 -32280 -23576 -30024
rect -16706 -30895 -16653 -30885
rect -16706 -31085 -16687 -30895
rect -16687 -31085 -16653 -30895
rect -16706 -31086 -16653 -31085
rect -16152 -30893 -16099 -30886
rect -16152 -31083 -16137 -30893
rect -16137 -31083 -16103 -30893
rect -16103 -31083 -16099 -30893
rect -16152 -31087 -16099 -31083
rect -15983 -31007 -15773 -30981
rect -15983 -31034 -15773 -31007
<< metal2 >>
rect -20400 3360 -9499 49600
rect -22348 422 -16669 423
rect -22350 -50 -16669 422
rect -22822 -1386 -16669 -50
rect -22342 -1388 -16669 -1386
rect -85199 -10677 -23576 -9757
rect -85199 -28067 -79389 -10677
rect -78189 -28067 -67389 -10677
rect -66189 -28067 -55389 -10677
rect -54189 -28067 -43389 -10677
rect -42189 -28067 -31389 -10677
rect -30189 -28067 -23576 -10677
rect -85199 -30024 -23576 -28067
rect -21900 -13290 -21160 -13280
rect -18340 -13418 -16669 -1388
rect -15440 -13300 -14700 -13290
rect -21900 -29420 -21160 -29410
rect -16566 -29414 -16506 -28852
rect -16682 -29474 -16506 -29414
rect -16462 -29415 -16402 -28852
rect -15440 -29410 -14700 -29400
rect -16682 -30389 -16622 -29474
rect -16462 -29475 -16262 -29415
rect -16322 -30310 -16262 -29475
rect -16322 -30363 -16100 -30310
rect -16707 -30444 -16622 -30389
rect -16707 -30590 -16654 -30444
rect -16153 -30590 -16100 -30363
rect -16706 -30885 -16653 -30590
rect -16706 -31094 -16653 -31086
rect -16152 -30886 -16099 -30590
rect -16152 -31095 -16099 -31087
rect -16024 -31034 -15983 -30981
rect -15773 -31034 -15765 -30981
rect -16024 -31378 -15987 -31034
rect -85199 -32290 -23576 -32280
rect -16682 -31438 -15987 -31378
rect -16682 -44204 -16622 -31438
<< via2 >>
rect -21900 -13300 -21160 -13290
rect -21900 -29400 -21500 -13300
rect -21500 -29400 -21160 -13300
rect -21900 -29410 -21160 -29400
rect -85199 -32280 -23576 -30024
rect -15440 -29400 -15100 -13300
rect -15100 -29400 -14700 -13300
<< metal3 >>
rect -89200 -4000 -79200 66802
rect -75200 56800 -9502 66800
rect -18400 43364 -9502 56800
rect -18400 3411 -9500 43364
rect -20400 1520 -9500 3411
rect -89200 -4576 -22388 -4000
rect -89200 -11276 -21135 -4576
rect -89200 -12561 -82816 -11276
rect -25932 -12561 -21135 -11276
rect -89200 -13290 -21135 -12561
rect -89200 -18044 -21900 -13290
rect -89200 -19329 -82559 -18044
rect -25675 -19329 -21900 -18044
rect -89200 -24000 -21900 -19329
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11471 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11471 -13300
rect -85209 -30024 -23566 -30019
rect -15464 -30024 -11471 -29400
rect -87200 -32280 -85199 -30024
rect -23576 -32280 -11471 -30024
rect -87200 -37148 -11471 -32280
rect -87200 -38433 -79646 -37148
rect -22762 -38433 -11471 -37148
rect -87200 -44000 -11471 -38433
<< via3 >>
rect -21900 -29410 -21160 -13290
rect -15440 -29400 -14700 -13300
rect -85199 -32280 -23576 -30024
<< metal4 >>
rect -89200 60593 -79200 66802
rect -89200 58735 -86553 60593
rect -81823 58735 -79200 60593
rect -89200 52593 -79200 58735
rect -75200 64072 -9502 66800
rect -75200 59258 -71351 64072
rect -69409 59258 -63351 64072
rect -61409 59258 -55351 64072
rect -53409 59258 -47351 64072
rect -45409 59258 -39351 64072
rect -37409 59258 -31351 64072
rect -29409 59258 -23351 64072
rect -21409 59258 -15351 64072
rect -13409 59258 -9502 64072
rect -75200 56800 -9502 59258
rect -89200 50735 -86553 52593
rect -81823 50735 -79200 52593
rect -89200 44593 -79200 50735
rect -89200 42735 -86553 44593
rect -81823 42735 -79200 44593
rect -89200 36593 -79200 42735
rect -89200 34735 -86553 36593
rect -81823 34735 -79200 36593
rect -89200 28593 -79200 34735
rect -89200 26735 -86553 28593
rect -81823 26735 -79200 28593
rect -89200 20593 -79200 26735
rect -89200 18735 -86553 20593
rect -81823 18735 -79200 20593
rect -89200 12593 -79200 18735
rect -89200 10735 -86553 12593
rect -81823 10735 -79200 12593
rect -89200 4593 -79200 10735
rect -89200 2735 -86553 4593
rect -81823 2735 -79200 4593
rect -18400 55488 -9502 56800
rect -18400 53376 -16710 55488
rect -12065 53376 -9502 55488
rect -18400 47488 -9502 53376
rect -18400 45376 -16710 47488
rect -12065 45376 -9502 47488
rect -18400 43364 -9502 45376
rect -18400 39488 -9500 43364
rect -18400 37376 -16710 39488
rect -12065 37376 -9500 39488
rect -18400 31488 -9500 37376
rect -18400 29376 -16710 31488
rect -12065 29376 -9500 31488
rect -18400 23488 -9500 29376
rect -18400 21376 -16710 23488
rect -12065 21376 -9500 23488
rect -18400 15488 -9500 21376
rect -18400 13376 -16710 15488
rect -12065 13376 -9500 15488
rect -18400 7488 -9500 13376
rect -18400 5376 -16710 7488
rect -12065 5376 -9500 7488
rect -18400 3411 -9500 5376
rect -89200 -3407 -79200 2735
rect -20400 1520 -9500 3411
rect -89200 -5265 -86553 -3407
rect -81823 -4000 -79200 -3407
rect -81823 -4576 -22388 -4000
rect -81823 -5265 -21135 -4576
rect -89200 -10417 -21135 -5265
rect -89200 -13288 -83681 -10417
rect -25493 -13288 -21135 -10417
rect -89200 -13290 -21135 -13288
rect -89200 -17342 -21900 -13290
rect -89200 -20213 -83343 -17342
rect -25155 -20213 -21900 -17342
rect -89200 -24000 -21900 -20213
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11471 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11471 -13300
rect -85200 -30024 -23575 -30023
rect -15464 -30024 -11471 -29400
rect -87200 -32280 -85199 -30024
rect -23576 -32280 -11471 -30024
rect -87200 -36344 -11471 -32280
rect -87200 -39215 -80725 -36344
rect -22537 -39215 -11471 -36344
rect -87200 -44000 -11471 -39215
<< via4 >>
rect -21900 -29410 -21160 -13290
rect -15440 -29400 -14700 -13300
rect -85199 -32280 -23576 -30024
<< metal5 >>
rect -89200 -4000 -79200 66802
rect -75200 56800 -9502 66800
rect -18400 43364 -9502 56800
rect -18400 3411 -9500 43364
rect -20400 1520 -9500 3411
rect -89200 -4576 -22388 -4000
rect -89200 -11276 -21135 -4576
rect -89200 -12561 -82816 -11276
rect -25932 -12561 -21135 -11276
rect -89200 -13290 -21135 -12561
rect -89200 -18044 -21900 -13290
rect -89200 -19329 -82559 -18044
rect -25675 -19329 -21900 -18044
rect -89200 -24000 -21900 -19329
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11471 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11471 -13300
rect -21924 -29434 -21136 -29433
rect -85223 -30024 -23552 -30000
rect -15464 -30024 -11471 -29400
rect -87200 -32280 -85199 -30024
rect -23576 -32280 -11471 -30024
rect -87200 -37148 -11471 -32280
rect -87200 -38433 -79646 -37148
rect -22762 -38433 -11471 -37148
rect -87200 -44000 -11471 -38433
use gate_drive  gate_drive_0
timestamp 1714671390
transform 0 -1 -17500 1 0 -20900
box -8928 -2874 8049 4445
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1714596710
transform -1 0 -22400 0 1 0
box -11346 -11351 64080 64140
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712845802
transform -1 0 -15249 0 1 -31230
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1712845802
transform -1 0 -16721 0 1 -31230
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712845802
transform -1 0 -15525 0 1 -31230
box -38 -48 222 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712845802
transform -1 0 -15709 0 1 -31230
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1712845802
transform -1 0 -16261 0 1 -31230
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712845802
transform -1 0 -15157 0 1 -31230
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1712845802
transform -1 0 -16169 0 1 -31230
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1712845802
transform -1 0 -16997 0 1 -31230
box -38 -48 130 592
<< labels >>
flabel metal5 -89200 66679 -79200 66802 5 FreeSans 8000 0 0 0 vdd_pwr
port 9 s
flabel metal5 -87200 -44000 -87179 -30024 1 FreeSans 8000 0 0 0 vss
port 10 n
flabel metal2 -16682 -44204 -16622 -44203 1 FreeSans 400 0 0 0 p_in
port 3 n
flabel metal5 -75200 65820 -9502 66800 1 FreeSans 8000 0 0 0 sw_node
port 7 n
flabel space -12049 -30733 -11477 -30254 0 FreeSans 4800 0 0 0 dvdd
port 11 nsew
flabel metal1 -12356 -12681 -11156 -11481 0 FreeSans 4800 0 0 0 dvss
port 6 nsew
<< end >>
