magic
tech sky130A
magscale 1 2
timestamp 1713985419
<< psubdiff >>
rect 3348 5238 3488 5296
rect 3348 4636 3382 5238
rect 3430 4636 3488 5238
rect 3348 4624 3488 4636
<< psubdiffcont >>
rect 3382 4636 3430 5238
<< locali >>
rect 2942 6450 3028 6470
rect 2942 6126 2952 6450
rect 3016 6126 3028 6450
rect 2942 6112 3028 6126
rect 1184 5502 1430 5506
rect -1418 5456 -974 5470
rect -1418 5412 -1404 5456
rect -990 5412 -974 5456
rect -1418 5398 -974 5412
rect -908 5456 -464 5470
rect -908 5412 -890 5456
rect -486 5412 -464 5456
rect -908 5398 -464 5412
rect 1184 5374 1202 5502
rect 1410 5374 1430 5502
rect 1184 5366 1430 5374
rect 3340 5238 3474 5286
rect -1190 4992 -702 5096
rect 3340 5074 3382 5238
rect 886 4922 3382 5074
rect -2108 4734 -1552 4762
rect -2108 4642 -2090 4734
rect -1570 4642 -1552 4734
rect -2108 4636 -1552 4642
rect 160 4712 3046 4722
rect 160 4638 166 4712
rect 3036 4638 3046 4712
rect 160 4632 3046 4638
rect 3340 4636 3382 4922
rect 3430 4636 3474 5238
<< viali >>
rect 2952 6126 3016 6450
rect -1404 5412 -990 5456
rect -890 5412 -486 5456
rect 1202 5374 1410 5502
rect -2090 4642 -1570 4734
rect 166 4638 3036 4712
<< metal1 >>
rect 896 6718 3020 6722
rect -1984 6234 410 6712
rect -1984 4780 -1518 6234
rect -1256 5802 -630 6234
rect -446 6054 -428 6148
rect -220 6054 -204 6148
rect -404 5470 -316 6054
rect -1418 5456 -974 5470
rect -1418 5412 -1404 5456
rect -990 5412 -974 5456
rect -1418 5398 -974 5412
rect -908 5456 -316 5470
rect -908 5412 -890 5456
rect -486 5412 -316 5456
rect -908 5398 -316 5412
rect -1418 5366 -1330 5398
rect -2218 4738 -1518 4780
rect -2218 4608 -2096 4738
rect -1588 4734 -1518 4738
rect -1570 4642 -1518 4734
rect -1588 4608 -1518 4642
rect -2218 4556 -1518 4608
rect -1420 4369 -1330 5366
rect -1248 5118 -462 5176
rect -1248 4942 -1198 5118
rect -516 4942 -462 5118
rect -1248 4890 -462 4942
rect -404 4352 -316 5398
rect -66 5802 410 6234
rect 558 6590 3020 6718
rect 558 6566 1128 6590
rect -66 4742 408 5802
rect 558 5182 816 6566
rect 2942 6460 3174 6470
rect 2942 6450 3090 6460
rect 2942 6126 2952 6450
rect 3016 6126 3090 6450
rect 2942 6122 3090 6126
rect 3158 6122 3174 6460
rect 2942 6112 3174 6122
rect 896 5760 3500 6004
rect 908 5694 2994 5710
rect 908 5642 948 5694
rect 2938 5642 2994 5694
rect 908 5630 2994 5642
rect 1184 5502 1430 5508
rect 1184 5374 1202 5502
rect 1410 5374 1430 5502
rect 1184 5366 1430 5374
rect 558 5176 1004 5182
rect 554 5082 3012 5176
rect 554 4958 928 5082
rect 2888 4958 3012 5082
rect 554 4890 3012 4958
rect 3218 4742 3500 5760
rect -66 4712 3500 4742
rect -66 4638 166 4712
rect -66 4602 226 4638
rect 3098 4602 3500 4712
rect -66 4530 3500 4602
rect -66 4528 408 4530
<< via1 >>
rect -428 6054 -220 6148
rect -2096 4734 -1588 4738
rect -2096 4642 -2090 4734
rect -2090 4642 -1588 4734
rect -2096 4608 -1588 4642
rect -1198 4942 -516 5118
rect 3090 6122 3158 6460
rect 948 5642 2938 5694
rect 1202 5374 1410 5502
rect 928 4958 2888 5082
rect 226 4638 3036 4712
rect 3036 4638 3098 4712
rect 226 4602 3098 4638
<< metal2 >>
rect 3082 6460 3168 6470
rect -446 6054 -428 6148
rect -220 6122 -204 6148
rect 3082 6122 3090 6460
rect 3158 6122 3168 6460
rect -220 6054 3174 6122
rect -2360 5918 -2050 5924
rect -2360 5694 2994 5918
rect -2360 5642 948 5694
rect 2938 5642 2994 5694
rect -2360 5614 2994 5642
rect 1184 5502 1430 5508
rect 1184 5494 1202 5502
rect -2370 5374 1202 5494
rect 1410 5374 1430 5502
rect -2370 5372 1430 5374
rect 1184 5366 1430 5372
rect -2384 5118 2944 5176
rect -2384 4942 -1198 5118
rect -516 5082 2944 5118
rect -516 4958 928 5082
rect 2888 4958 2944 5082
rect -516 4942 2944 4958
rect -2384 4890 2944 4942
rect -2394 4738 3498 4814
rect -2394 4608 -2096 4738
rect -1588 4712 3498 4738
rect -1588 4608 226 4712
rect -2394 4602 226 4608
rect 3098 4602 3498 4712
rect -2394 4506 3498 4602
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform -1 0 -704 0 1 5089
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1712845802
transform 1 0 896 0 1 5065
box -66 -43 2178 1671
<< labels >>
flabel metal1 -404 4352 -316 4432 0 FreeSans 560 0 0 0 out3v3
port 9 nsew
flabel metal1 -1420 4369 -1330 4459 0 FreeSans 560 0 0 0 outb3v3
port 10 nsew
flabel metal2 -2370 5372 -2048 5494 0 FreeSans 560 0 0 0 in1v8
port 1 nsew
flabel metal2 -2394 4506 -2106 4814 0 FreeSans 560 0 0 0 avdd
port 8 nsew
flabel metal2 -2384 4890 -2052 5176 0 FreeSans 560 0 0 0 dvss
port 0 nsew
flabel metal2 -2360 5614 -2050 5924 0 FreeSans 560 0 0 0 dvdd
port 2 nsew
<< end >>
