magic
tech sky130A
magscale 1 2
timestamp 1715098825
<< isosubstrate >>
rect 800 649276 282072 704800
rect 800 574016 170892 649276
rect 246180 645694 282072 649276
rect 246180 638530 247856 645694
rect 264692 638530 282072 645694
rect 246180 574016 282072 638530
rect 800 559258 282072 574016
rect 800 540902 170890 559258
rect 800 482300 4146 540902
rect 20326 482300 22616 484688
rect 26908 483998 170890 540902
rect 246178 555704 282072 559258
rect 246178 548540 247840 555704
rect 264676 548540 282072 555704
rect 246178 483998 282072 548540
rect 26908 482300 282072 483998
rect 800 469256 282072 482300
rect 800 466376 170874 469256
rect 800 462114 5296 466376
rect 8524 465452 170874 466376
rect 10130 462114 170874 465452
rect 800 461174 170874 462114
rect 800 456916 5300 461174
rect 10130 457826 170874 461174
rect 8528 456916 170874 457826
rect 800 432550 170874 456916
rect 800 432540 7198 432550
rect 800 430948 2902 432540
rect 800 427704 1984 430948
rect 6244 427710 7198 432540
rect 10526 430948 170874 432550
rect 11464 427710 170874 430948
rect 6244 427704 170874 427710
rect 800 393996 170874 427704
rect 246162 465704 282072 469256
rect 246162 458540 247856 465704
rect 264692 458540 282072 465704
rect 246162 393996 282072 458540
rect 800 384936 282072 393996
rect 800 381694 2976 384936
rect 800 380098 3876 381694
rect 7228 380098 282072 384936
rect 800 379268 282072 380098
rect 800 358830 170890 379268
rect 800 353890 21092 358830
rect 59660 353890 170890 358830
rect 800 349788 16880 353890
rect 59682 351310 170890 353890
rect 61754 349788 170890 351310
rect 800 344226 14972 349788
rect 800 339908 2744 344226
rect 6054 343300 14972 344226
rect 7638 339908 14972 343300
rect 800 339034 14972 339908
rect 800 334738 2744 339034
rect 7626 335612 14972 339034
rect 6012 334738 14972 335612
rect 800 317808 14972 334738
rect 61776 317808 170890 349788
rect 800 304008 170890 317808
rect 246178 375698 282072 379268
rect 246178 368534 247848 375698
rect 264684 368534 282072 375698
rect 246178 304008 282072 368534
rect 800 301028 282072 304008
rect 800 296748 3188 301028
rect 6458 300100 282072 301028
rect 8052 299748 282072 300100
rect 8052 299746 40550 299748
rect 8052 296748 17528 299746
rect 800 295862 17528 296748
rect 800 291576 3188 295862
rect 6454 295858 17528 295862
rect 8058 292444 17528 295858
rect 6454 291576 17528 292444
rect 800 220520 17528 291576
rect 25548 220522 40550 299746
rect 48570 289258 282072 299748
rect 48570 220522 170876 289258
rect 25548 220520 170876 220522
rect 800 213998 170876 220520
rect 246164 285708 282072 289258
rect 246164 278544 247854 285708
rect 264690 278544 282072 285708
rect 246164 213998 282072 278544
rect 800 199262 282072 213998
rect 800 124002 170874 199262
rect 246162 195688 282072 199262
rect 246162 188524 247856 195688
rect 264692 188524 282072 195688
rect 246162 124002 282072 188524
rect 800 110748 282072 124002
rect 800 98494 12730 110748
rect 20322 109264 282072 110748
rect 20322 108978 170898 109264
rect 20322 98494 23266 108978
rect 800 96848 23266 98494
rect 800 91122 12154 96848
rect 17284 93570 23266 96848
rect 33188 98044 33974 108978
rect 36742 98044 170898 108978
rect 33188 93570 170898 98044
rect 17284 91122 170898 93570
rect 800 56598 170898 91122
rect 800 56552 38702 56598
rect 800 49666 32896 56552
rect 37640 49666 38702 56552
rect 800 43934 38702 49666
rect 800 39616 3350 43934
rect 6684 43006 38702 43934
rect 8278 42834 38702 43006
rect 59846 56584 170898 56598
rect 59846 42834 60870 56584
rect 8278 42794 60870 42834
rect 79976 42794 170898 56584
rect 8278 39616 170898 42794
rect 800 38778 170898 39616
rect 800 38772 6592 38778
rect 800 34410 3368 38772
rect 8278 35308 170898 38778
rect 6684 34410 170898 35308
rect 800 34004 170898 34410
rect 246186 105702 282072 109264
rect 246186 98538 247854 105702
rect 264690 98538 282072 105702
rect 246186 34004 282072 98538
rect 800 800 282072 34004
rect 282270 649226 584800 704800
rect 282270 645710 340600 649226
rect 282270 638542 322104 645710
rect 338944 638542 340600 645710
rect 282270 574000 340600 638542
rect 415916 594390 584800 649226
rect 415916 574000 521090 594390
rect 545696 592364 584800 594390
rect 545696 586816 547194 592364
rect 545696 585994 550746 586816
rect 282270 572486 521090 574000
rect 549924 575980 550746 585994
rect 563724 586732 584800 592364
rect 563724 586726 582732 586732
rect 563724 581838 579398 586726
rect 583718 583472 584800 586732
rect 582806 581838 584800 583472
rect 563724 575980 584800 581838
rect 549924 572486 584800 575980
rect 282270 559238 584800 572486
rect 282270 555706 340608 559238
rect 282270 548538 322084 555706
rect 338924 548538 340608 555706
rect 282270 484012 340608 548538
rect 415924 497246 584800 559238
rect 415924 497240 582282 497246
rect 415924 492398 579018 497240
rect 583298 494004 584800 497246
rect 582400 492398 584800 494004
rect 415924 484012 584800 492398
rect 282270 469234 584800 484012
rect 282270 465698 340618 469234
rect 282270 458530 322106 465698
rect 338946 458530 340618 465698
rect 282270 394008 340618 458530
rect 415934 436354 584800 469234
rect 415934 436140 569998 436354
rect 415934 419394 562584 436140
rect 568904 419394 569998 436140
rect 415934 417294 569998 419394
rect 415934 412542 561784 417294
rect 567586 412542 569998 417294
rect 415934 412328 569998 412542
rect 582208 412328 584800 436354
rect 415934 394008 584800 412328
rect 282270 379236 584800 394008
rect 282270 375710 340602 379236
rect 282270 368542 322096 375710
rect 338936 368542 340602 375710
rect 282270 304010 340602 368542
rect 415918 365628 584800 379236
rect 415918 364726 580102 365628
rect 583378 364726 584800 365628
rect 415918 361338 578554 364726
rect 583392 361338 584800 364726
rect 415918 360400 584800 361338
rect 415918 357042 578554 360400
rect 415918 356156 580154 357042
rect 583370 356156 584800 360400
rect 415918 316822 584800 356156
rect 415918 316814 576290 316822
rect 415918 311996 573044 316814
rect 577280 313568 584800 316822
rect 576386 311996 584800 313568
rect 415918 304010 584800 311996
rect 282270 294538 584800 304010
rect 282270 289226 517066 294538
rect 536592 294504 584800 294538
rect 282270 285708 340594 289226
rect 282270 282484 322090 285708
rect 282270 32326 289370 282484
rect 297538 278540 322090 282484
rect 338930 278540 340594 285708
rect 297538 214000 340594 278540
rect 415910 271446 517066 289226
rect 555802 281262 584800 294504
rect 551352 280556 584800 281262
rect 530908 271446 536380 275400
rect 415910 270598 536380 271446
rect 415910 267456 517736 270598
rect 520808 270564 536380 270598
rect 520808 267456 525046 270564
rect 415910 265972 525046 267456
rect 531648 265972 536380 270564
rect 415910 252766 536380 265972
rect 551352 252766 552226 280556
rect 415910 251940 552226 252766
rect 557178 272368 584800 280556
rect 557178 272360 582698 272368
rect 557178 267508 579420 272360
rect 583676 269120 584800 272368
rect 582780 267508 584800 269120
rect 557178 251940 584800 267508
rect 415910 214000 584800 251940
rect 297538 199234 584800 214000
rect 297538 195712 340602 199234
rect 297538 188536 322092 195712
rect 338914 188536 340602 195712
rect 297538 124008 340602 188536
rect 415918 177814 584800 199234
rect 415918 154626 522854 177814
rect 533892 177754 584800 177814
rect 533892 154626 539306 158536
rect 415918 153662 539306 154626
rect 415918 150534 523546 153662
rect 526524 153632 539306 153662
rect 526524 150534 527486 153632
rect 415918 149752 527486 150534
rect 534494 149752 539306 153632
rect 415918 136068 539306 149752
rect 550826 136068 584800 177754
rect 415918 124008 584800 136068
rect 297538 109240 584800 124008
rect 297538 105714 340592 109240
rect 297538 98538 322098 105714
rect 338920 98538 340592 105714
rect 297538 34014 340592 98538
rect 415908 88878 584800 109240
rect 415908 65842 517478 88878
rect 556020 75770 584800 88878
rect 551670 74870 584800 75770
rect 531304 65842 536734 69862
rect 415908 64972 536734 65842
rect 415908 61942 518078 64972
rect 521166 64942 536734 64972
rect 521166 61942 522216 64942
rect 415908 60444 522216 61942
rect 531904 60444 536734 64942
rect 415908 47276 536734 60444
rect 551670 47366 552420 74870
rect 557518 47366 584800 74870
rect 551670 47276 584800 47366
rect 415908 34014 584800 47276
rect 297538 32326 584800 34014
rect 282270 800 584800 32326
<< metal1 >>
rect 263426 654713 265741 654863
rect 263426 653984 263662 654713
rect 265591 653984 265741 654713
rect 263426 653791 265741 653984
rect 321050 654704 323365 654854
rect 321050 653975 321200 654704
rect 323129 653975 323365 654704
rect 245574 653106 247889 653256
rect 245574 652377 245788 653106
rect 247717 652377 247889 653106
rect 245574 652184 247889 652377
rect 246275 651795 247829 652184
rect 246277 649354 247829 651795
rect 246276 649161 247829 649354
rect 265195 648781 265674 653791
rect 321050 653782 323365 653975
rect 321117 648486 321596 653782
rect 338902 653097 341217 653247
rect 338902 652368 339074 653097
rect 341003 652368 341217 653097
rect 338902 652175 341217 652368
rect 338962 649156 340516 652175
rect 513415 609778 520733 610315
rect 508780 594670 510602 595116
rect 513415 595070 513911 609778
rect 513414 594741 513911 595070
rect 513415 593259 513911 594741
rect 520276 594202 520733 609778
rect 556287 601770 560183 602040
rect 520276 593259 521512 594202
rect 556287 593934 556508 601770
rect 560007 593934 560183 601770
rect 556287 593698 560183 593934
rect 513415 592789 521512 593259
rect 573463 586727 574467 586813
rect 573463 585613 573573 586727
rect 574366 586445 574467 586727
rect 574366 586209 579592 586445
rect 574366 585613 574467 586209
rect 573463 585534 574467 585613
rect 567699 584944 579640 585047
rect 567699 580597 567802 584944
rect 583830 584564 584262 584602
rect 583830 584468 583874 584564
rect 583634 584326 583874 584468
rect 583830 584260 583874 584326
rect 584212 584260 584262 584564
rect 583830 584232 584262 584260
rect 577087 584173 577726 584230
rect 577087 584083 577145 584173
rect 577085 583814 577145 584083
rect 577087 583409 577145 583814
rect 577661 584083 577726 584173
rect 577661 583814 579591 584083
rect 577661 583409 577726 583814
rect 577087 583360 577726 583409
rect 578078 581725 579692 581749
rect 578078 581498 578165 581725
rect 579312 581498 579692 581725
rect 578078 581465 579692 581498
rect 567629 580543 567862 580597
rect 567629 579827 567667 580543
rect 567829 579827 567862 580543
rect 567629 579773 567862 579827
rect 510422 576926 518844 577547
rect 510422 570179 510907 576926
rect 518330 574012 518844 576926
rect 518330 572711 521727 574012
rect 556374 572886 560268 573078
rect 518330 570179 518844 572711
rect 510422 569612 518844 570179
rect 263426 564713 265741 564863
rect 263426 563984 263662 564713
rect 265591 563984 265741 564713
rect 263426 563791 265741 563984
rect 321050 564704 323365 564854
rect 321050 563975 321200 564704
rect 323129 563975 323365 564704
rect 245574 563106 247889 563256
rect 245574 562377 245788 563106
rect 247717 562377 247889 563106
rect 245574 562184 247889 562377
rect 246275 561795 247829 562184
rect 246277 559354 247829 561795
rect 246276 559161 247829 559354
rect 265195 558781 265674 563791
rect 321050 563782 323365 563975
rect 321117 558486 321596 563782
rect 338902 563097 341217 563247
rect 338902 562368 339074 563097
rect 341003 562368 341217 563097
rect 556374 563187 556611 572886
rect 560065 563187 560268 572886
rect 556374 562979 560268 563187
rect 338902 562175 341217 562368
rect 338962 559156 340516 562175
rect 575990 498421 576687 498523
rect 575990 496743 576075 498421
rect 576616 496994 576687 498421
rect 576616 496767 579231 496994
rect 576616 496743 576687 496767
rect 575990 496650 576687 496743
rect 574914 496291 575907 496393
rect 574914 495447 575013 496291
rect 575808 495668 575907 496291
rect 575808 495460 579161 495668
rect 575808 495447 575907 495460
rect 574914 495358 575907 495447
rect 583438 495102 584234 495148
rect 583438 495044 583490 495102
rect 576700 494849 577862 494922
rect 583226 494920 583490 495044
rect 576700 493993 576790 494849
rect 577757 494660 577862 494849
rect 583438 494882 583490 494920
rect 584168 494882 584234 495102
rect 583438 494838 584234 494882
rect 577757 494395 579163 494660
rect 577757 493993 577862 494395
rect 576700 493929 577862 493993
rect 578266 492276 579461 492320
rect 578266 492070 578317 492276
rect 579412 492070 579461 492276
rect 578266 492032 579461 492070
rect 4613 475393 6213 482370
rect 20479 480490 20752 482778
rect 20445 480450 20812 480490
rect 20445 479565 20480 480450
rect 20783 479565 20812 480450
rect 20445 479522 20812 479565
rect 21251 476758 21407 482669
rect 22022 481278 22295 482788
rect 21973 481235 22340 481278
rect 21973 480350 22005 481235
rect 22308 480350 22340 481235
rect 21973 480310 22340 480350
rect 263426 477313 265741 477463
rect 21251 476743 21774 476758
rect 21251 476599 21268 476743
rect 21751 476599 21774 476743
rect 21251 476583 21774 476599
rect 263426 476584 263662 477313
rect 265591 476584 265741 477313
rect 263426 476391 265741 476584
rect 4613 470506 4728 475393
rect 6108 470506 6213 475393
rect 245574 473106 247889 473256
rect 245574 472377 245788 473106
rect 247717 472377 247889 473106
rect 245574 472184 247889 472377
rect 246275 471795 247829 472184
rect 4613 470387 6213 470506
rect 4745 470220 6027 470387
rect 246277 469354 247829 471795
rect 246276 469161 247829 469354
rect 265195 468781 265674 476391
rect 321050 474704 323365 474854
rect 321050 473975 321200 474704
rect 323129 473975 323365 474704
rect 321050 473782 323365 473975
rect 321117 468486 321596 473782
rect 338902 473097 341217 473247
rect 338902 472368 339074 473097
rect 341003 472368 341217 473097
rect 338902 472175 341217 472368
rect 338962 469156 340516 472175
rect 7456 468312 7723 468354
rect 7456 467721 7486 468312
rect 7690 467721 7723 468312
rect 7456 467681 7723 467721
rect 7468 466529 7714 467681
rect 7466 461984 8347 462028
rect 2167 461759 5322 461778
rect 2167 461534 2194 461759
rect 3030 461534 5322 461759
rect 2167 461516 5322 461534
rect 7466 461352 7523 461984
rect 8290 461352 8347 461984
rect 7466 461302 8347 461352
rect 7483 455643 7697 456871
rect 7345 455429 7697 455643
rect 7345 443441 7559 455429
rect 9023 448336 10305 448514
rect 9023 446702 9147 448336
rect 10216 446702 10305 448336
rect 9023 444149 10305 446702
rect 7345 443227 9245 443441
rect 6462 439485 6743 439503
rect 6462 438897 6476 439485
rect 6728 439467 6743 439485
rect 6728 439345 9627 439467
rect 6728 438897 6743 439345
rect 6462 438880 6743 438897
rect 7368 439022 7592 439029
rect 7368 439002 9597 439022
rect 7368 438204 7391 439002
rect 7570 438909 9597 439002
rect 7570 438204 7592 438909
rect 7368 438178 7592 438204
rect 7959 438229 9673 438469
rect 1703 435904 2427 435927
rect 1703 435716 1738 435904
rect 2398 435716 2427 435904
rect 1703 435690 2427 435716
rect 1747 429872 1993 435690
rect 7959 435555 8199 438229
rect 13208 437642 14598 437666
rect 13208 437442 13238 437642
rect 14564 437442 14598 437642
rect 13208 437416 14598 437442
rect 7959 435315 11729 435555
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 6302 429814 7162 429877
rect 11489 429872 11729 435315
rect 4484 426541 4759 426576
rect 4484 425868 4522 426541
rect 4717 426147 4759 426541
rect 6577 426147 6839 427726
rect 4717 425885 6839 426147
rect 4717 425868 4759 425885
rect 4484 425830 4759 425868
rect 8087 384757 9234 384793
rect 8087 384667 8126 384757
rect 7065 384475 8126 384667
rect 9182 384475 9234 384757
rect 7065 384444 9234 384475
rect 8087 384441 9234 384444
rect 263426 384713 265741 384863
rect 263426 383984 263662 384713
rect 265591 383984 265741 384713
rect 263426 383791 265741 383984
rect 321050 384704 323365 384854
rect 321050 383975 321200 384704
rect 323129 383975 323365 384704
rect 8490 383334 9178 383354
rect 7139 383290 9178 383334
rect 7139 383132 8553 383290
rect 8490 382858 8553 383132
rect 9115 382858 9178 383290
rect 1694 382780 2576 382812
rect 8490 382807 9178 382858
rect 245574 383106 247889 383256
rect 1694 382608 1730 382780
rect 2548 382718 2576 382780
rect 2548 382608 3102 382718
rect 1694 382598 3102 382608
rect 1694 382578 2576 382598
rect 245574 382377 245788 383106
rect 247717 382377 247889 383106
rect 8167 382336 9436 382347
rect 7090 382289 9436 382336
rect 7090 382065 8241 382289
rect 8167 381897 8241 382065
rect 9368 381897 9436 382289
rect 245574 382184 247889 382377
rect 8167 381846 9436 381897
rect 246275 381795 247829 382184
rect 7571 380014 9262 380019
rect 6839 379992 9262 380014
rect 6839 379740 7617 379992
rect 9223 379740 9262 379992
rect 6839 379709 9262 379740
rect 6839 379706 8545 379709
rect 246277 379254 247829 381795
rect 265195 378844 265674 383791
rect 321050 383782 323365 383975
rect 321117 378486 321596 383782
rect 338902 383097 341217 383247
rect 338902 382368 339074 383097
rect 341003 382368 341217 383097
rect 338902 382175 341217 382368
rect 338962 379156 340516 382175
rect 580981 367266 581227 367315
rect 580981 365564 581227 366286
rect 580109 361187 581287 361243
rect 580109 360563 580208 361187
rect 581211 360563 581287 361187
rect 583575 361027 584320 361051
rect 583575 360769 583603 361027
rect 584293 360769 584320 361027
rect 583575 360746 584320 360769
rect 580109 360507 581287 360563
rect 59776 359034 60384 359062
rect 59776 358268 59802 359034
rect 60356 358268 60384 359034
rect 59776 358236 60384 358268
rect 580987 355293 581227 355892
rect 580987 354384 581001 355293
rect 580987 354365 581227 354384
rect 4957 344582 5920 344626
rect 4957 344467 4993 344582
rect 5879 344467 5920 344582
rect 4957 344428 5920 344467
rect 4935 339653 6035 339688
rect 1528 339574 2590 339613
rect 1528 339376 1564 339574
rect 2527 339376 2590 339574
rect 1528 339348 2590 339376
rect 4935 339220 4983 339653
rect 5982 339220 6035 339653
rect 4935 339168 6035 339220
rect 4943 334449 5832 334464
rect 4943 334263 4974 334449
rect 5809 334263 5832 334449
rect 4943 334244 5832 334263
rect 567090 316809 568186 316873
rect 567090 315844 567177 316809
rect 568123 316556 568186 316809
rect 568123 316328 573167 316556
rect 568123 315844 568186 316328
rect 567090 315777 568186 315844
rect 569251 315568 570067 315681
rect 569251 314111 569330 315568
rect 569965 315211 570067 315568
rect 569965 315013 573167 315211
rect 569965 314111 570067 315013
rect 582578 314662 583714 314710
rect 582578 314574 582644 314662
rect 577210 314468 582644 314574
rect 569251 313992 570067 314111
rect 571015 314309 572629 314379
rect 571015 313895 571103 314309
rect 572537 314215 572629 314309
rect 582578 314328 582644 314468
rect 583666 314328 583714 314662
rect 582578 314280 583714 314328
rect 572537 313936 573194 314215
rect 572537 313895 572629 313936
rect 571015 313812 572629 313895
rect 571839 311837 573546 311870
rect 571839 311649 571913 311837
rect 573518 311649 573546 311837
rect 571839 311590 573546 311649
rect 5372 301415 6335 301432
rect 5372 301251 5395 301415
rect 6315 301251 6335 301415
rect 5372 301234 6335 301251
rect 5194 296534 6467 296612
rect 1917 296389 2979 296430
rect 1917 296191 1959 296389
rect 2922 296191 2979 296389
rect 1917 296165 2979 296191
rect 5194 296044 5290 296534
rect 6335 296044 6467 296534
rect 5194 295966 6467 296044
rect 338902 295097 341217 295247
rect 263426 294713 265741 294863
rect 263426 293984 263662 294713
rect 265591 293984 265741 294713
rect 338902 294368 339074 295097
rect 341003 294368 341217 295097
rect 338902 294175 341217 294368
rect 263426 293791 265741 293984
rect 245574 293106 247889 293256
rect 245574 292377 245788 293106
rect 247717 292377 247889 293106
rect 245574 292184 247889 292377
rect 246275 291795 247829 292184
rect 5372 291271 6070 291289
rect 5372 291105 5396 291271
rect 6049 291105 6070 291271
rect 5372 291088 6070 291105
rect 246277 289228 247829 291795
rect 265195 288790 265674 293791
rect 321062 292916 323377 293065
rect 321062 292187 321212 292916
rect 323141 292187 323377 292916
rect 321062 291994 323377 292187
rect 321117 291992 321608 291994
rect 321117 288486 321596 291992
rect 338962 289156 340516 294175
rect 11135 286547 11237 286561
rect 11135 286443 11151 286547
rect 9757 286355 11151 286443
rect 11135 286351 11151 286355
rect 11227 286351 11237 286547
rect 11135 286333 11237 286351
rect 10965 285546 11073 285560
rect 10965 285429 10980 285546
rect 9738 285344 10980 285429
rect 11060 285429 11073 285546
rect 11060 285344 11084 285429
rect 9738 285339 11084 285344
rect 10965 285328 11073 285339
rect 578786 272103 579326 272134
rect 578786 272101 579726 272103
rect 578786 271811 578848 272101
rect 579290 271871 579726 272101
rect 579290 271811 579326 271871
rect 578786 271784 579326 271811
rect 578267 270783 579168 270845
rect 578267 270535 578316 270783
rect 579119 270764 579168 270783
rect 579119 270565 579524 270764
rect 579119 270535 579168 270565
rect 578267 270495 579168 270535
rect 583850 270272 584276 270316
rect 583850 270152 583912 270272
rect 583616 270016 583912 270152
rect 583850 269860 583912 270016
rect 584220 269860 584276 270272
rect 578265 269759 579153 269826
rect 583850 269812 584276 269860
rect 578262 269758 579541 269759
rect 578262 269501 578330 269758
rect 578265 269456 578330 269501
rect 579103 269501 579541 269758
rect 579103 269456 579153 269501
rect 578265 269412 579153 269456
rect 579005 267379 579830 267422
rect 579005 267185 579061 267379
rect 579777 267185 579830 267379
rect 579005 267142 579830 267185
rect 263426 204713 265741 204863
rect 263426 203984 263662 204713
rect 265591 203984 265741 204713
rect 263426 203791 265741 203984
rect 321050 204704 323365 204854
rect 321050 203975 321200 204704
rect 323129 203975 323365 204704
rect 245574 203106 247889 203256
rect 245574 202377 245788 203106
rect 247717 202377 247889 203106
rect 245574 202184 247889 202377
rect 246275 201795 247829 202184
rect 246277 199354 247829 201795
rect 246276 199161 247829 199354
rect 265195 198781 265674 203791
rect 321050 203782 323365 203975
rect 321117 198486 321596 203782
rect 338902 203097 341217 203247
rect 338902 202368 339074 203097
rect 341003 202368 341217 203097
rect 338902 202175 341217 202368
rect 338962 199156 340516 202175
rect 263426 114713 265741 114863
rect 263426 113984 263662 114713
rect 265591 113984 265741 114713
rect 263426 113791 265741 113984
rect 321050 114704 323365 114854
rect 321050 113975 321200 114704
rect 323129 113975 323365 114704
rect 245574 113106 247889 113256
rect 245574 112377 245788 113106
rect 247717 112377 247889 113106
rect 245574 112184 247889 112377
rect 246275 111795 247829 112184
rect 246277 109161 247829 111795
rect 265195 108914 265674 113791
rect 321050 113782 323365 113975
rect 321117 108452 321596 113782
rect 338902 113097 341217 113247
rect 338902 112368 339074 113097
rect 341003 112368 341217 113097
rect 338902 112175 341217 112368
rect 338962 109163 340516 112175
rect 265195 107747 265674 107947
rect 5595 44369 5844 44392
rect 5595 44084 5614 44369
rect 5821 44084 5844 44369
rect 5595 44063 5844 44084
rect 1456 39496 1714 39528
rect 1456 38894 1484 39496
rect 1684 39240 1714 39496
rect 5652 39422 6511 39493
rect 1684 39086 3448 39240
rect 1684 38894 1714 39086
rect 1456 38866 1714 38894
rect 5652 38923 5712 39422
rect 6434 38923 6511 39422
rect 5652 38883 6511 38923
rect 5623 34064 5817 34342
rect 5623 33870 7527 34064
rect 7333 28442 7527 33870
rect 290311 30949 290511 32541
rect 290073 30905 290992 30949
rect 290073 30361 290122 30905
rect 290933 30361 290992 30905
rect 290073 30317 290992 30361
rect 7204 28409 7656 28442
rect 7204 27214 7258 28409
rect 7592 27214 7656 28409
rect 7204 27149 7656 27214
<< via1 >>
rect 263662 653984 265591 654713
rect 321200 653975 323129 654704
rect 245788 652377 247717 653106
rect 339074 652368 341003 653097
rect 513911 593259 520276 609778
rect 556508 593934 560007 601770
rect 573573 585613 574366 586727
rect 583874 584260 584212 584564
rect 577145 583409 577661 584173
rect 578165 581498 579312 581725
rect 567667 579827 567829 580543
rect 510907 570179 518330 576926
rect 263662 563984 265591 564713
rect 321200 563975 323129 564704
rect 245788 562377 247717 563106
rect 339074 562368 341003 563097
rect 556611 563187 560065 572886
rect 25460 486521 26354 500270
rect 576075 496743 576616 498421
rect 575013 495447 575808 496291
rect 576790 493993 577757 494849
rect 583490 494882 584168 495102
rect 578317 492070 579412 492276
rect 20480 479565 20783 480450
rect 22005 480350 22308 481235
rect 21268 476599 21751 476743
rect 263662 476584 265591 477313
rect 4728 470506 6108 475393
rect 245788 472377 247717 473106
rect 321200 473975 323129 474704
rect 339074 472368 341003 473097
rect 7486 467721 7690 468312
rect 2194 461534 3030 461759
rect 7523 461352 8290 461984
rect 9147 446702 10216 448336
rect 6476 438897 6728 439485
rect 7391 438204 7570 439002
rect 1738 435716 2398 435904
rect 13238 437442 14564 437642
rect 6378 429877 7086 430832
rect 4522 425868 4717 426541
rect 8126 384475 9182 384757
rect 263662 383984 265591 384713
rect 321200 383975 323129 384704
rect 8553 382858 9115 383290
rect 1730 382608 2548 382780
rect 245788 382377 247717 383106
rect 8241 381897 9368 382289
rect 7617 379740 9223 379992
rect 339074 382368 341003 383097
rect 580981 366286 581227 367266
rect 580208 360563 581211 361187
rect 583603 360769 584293 361027
rect 59802 358268 60356 359034
rect 581001 354384 581227 355293
rect 4993 344467 5879 344582
rect 1564 339376 2527 339574
rect 4983 339220 5982 339653
rect 4974 334263 5809 334449
rect 567177 315844 568123 316809
rect 569330 314111 569965 315568
rect 571103 313895 572537 314309
rect 582644 314328 583666 314662
rect 571913 311649 573518 311837
rect 5395 301251 6315 301415
rect 1959 296191 2922 296389
rect 5290 296044 6335 296534
rect 263662 293984 265591 294713
rect 339074 294368 341003 295097
rect 245788 292377 247717 293106
rect 5396 291105 6049 291271
rect 321212 292187 323141 292916
rect 11151 286351 11227 286547
rect 10980 285344 11060 285546
rect 578848 271811 579290 272101
rect 578316 270535 579119 270783
rect 583912 269860 584220 270272
rect 578330 269456 579103 269758
rect 579061 267185 579777 267379
rect 263662 203984 265591 204713
rect 321200 203975 323129 204704
rect 245788 202377 247717 203106
rect 339074 202368 341003 203097
rect 263662 113984 265591 114713
rect 321200 113975 323129 114704
rect 245788 112377 247717 113106
rect 339074 112368 341003 113097
rect 5614 44084 5821 44369
rect 1484 38894 1684 39496
rect 5712 38923 6434 39422
rect 290122 30361 290933 30905
rect 7258 27214 7592 28409
<< metal2 >>
rect 263426 654713 265741 654863
rect 263426 653984 263662 654713
rect 265591 653984 265741 654713
rect 263426 653791 265741 653984
rect 321050 654704 323365 654854
rect 321050 653975 321200 654704
rect 323129 653975 323365 654704
rect 321050 653782 323365 653975
rect 245574 653106 247889 653256
rect 245574 652377 245788 653106
rect 247717 652377 247889 653106
rect 245574 652184 247889 652377
rect 338902 653097 341217 653247
rect 338902 652368 339074 653097
rect 341003 652368 341217 653097
rect 338902 652175 341217 652368
rect 279035 643726 282767 643786
rect 263426 564713 265741 564863
rect 263426 563984 263662 564713
rect 265591 563984 265741 564713
rect 263426 563791 265741 563984
rect 245574 563106 247889 563256
rect 245574 562377 245788 563106
rect 247717 562377 247889 563106
rect 245574 562184 247889 562377
rect 279035 553726 282487 553786
rect 25311 500270 26552 500469
rect 25311 492593 25460 500270
rect 25262 486521 25460 492593
rect 26354 492593 26552 500270
rect 26354 492430 38581 492593
rect 26354 486659 28395 492430
rect 38334 486659 38581 492430
rect 26354 486521 38581 486659
rect 25262 486422 38581 486521
rect 25311 486372 26552 486422
rect 4420 475393 12415 475493
rect 4420 470506 4728 475393
rect 6108 470506 6256 475393
rect 4420 470365 6256 470506
rect 12269 470365 12415 475393
rect 4420 470219 12415 470365
rect 15695 469792 15851 482422
rect 15621 469755 15920 469792
rect 2247 469256 2511 469276
rect 2247 468578 2262 469256
rect 2494 468578 2511 469256
rect 7459 469236 8334 469270
rect 7459 469100 7494 469236
rect 8300 469100 8334 469236
rect 7459 469073 8334 469100
rect 15621 469083 15660 469755
rect 15889 469083 15920 469755
rect 2247 468557 2511 468578
rect 2268 461777 2475 468557
rect 7505 468354 7690 469073
rect 15621 469053 15920 469083
rect 7456 468312 7723 468354
rect 7456 467721 7486 468312
rect 7690 467721 7723 468312
rect 7456 467681 7723 467721
rect 16967 467330 17123 482466
rect 18306 479594 18658 482471
rect 21973 481235 22340 481278
rect 20445 480450 20812 480490
rect 18196 479537 18710 479594
rect 18196 478121 18241 479537
rect 18645 478121 18710 479537
rect 20445 479565 20480 480450
rect 20783 479975 20812 480450
rect 21973 480350 22005 481235
rect 22308 480747 22340 481235
rect 136829 481050 140840 481122
rect 136829 480747 136929 481050
rect 22308 480414 136929 480747
rect 140755 480747 140840 481050
rect 140755 480414 140936 480747
rect 22308 480350 140936 480414
rect 21973 480346 140936 480350
rect 21973 480310 22340 480346
rect 128830 479975 132831 479982
rect 20783 479922 140936 479975
rect 20783 479574 128886 479922
rect 20783 479565 20812 479574
rect 20445 479522 20812 479565
rect 128830 479271 128886 479574
rect 132750 479574 140936 479922
rect 132750 479271 132831 479574
rect 128830 479211 132831 479271
rect 18196 478064 18710 478121
rect 263426 477313 265741 477463
rect 21251 476743 21774 476758
rect 21251 476599 21268 476743
rect 21751 476733 21774 476743
rect 21751 476633 142568 476733
rect 21751 476599 21774 476633
rect 21251 476583 21774 476599
rect 4524 467174 17123 467330
rect 2166 461759 3055 461777
rect 2166 461534 2194 461759
rect 3030 461534 3055 461759
rect 2166 461517 3055 461534
rect 2268 461516 2475 461517
rect 1703 435904 2427 435927
rect 1703 435716 1738 435904
rect 2398 435889 2427 435904
rect 4524 435889 4680 467174
rect 7466 461984 8347 462028
rect 7466 461352 7523 461984
rect 8290 461352 8347 461984
rect 7466 461302 8347 461352
rect 5382 456631 5786 456990
rect 5343 456528 6129 456631
rect 5343 455115 5436 456528
rect 6072 455115 6129 456528
rect 10238 456434 10524 458058
rect 10720 457049 10842 458191
rect 10962 458053 140941 458106
rect 10962 457796 136913 458053
rect 136832 457377 136913 457796
rect 140759 457796 140941 458053
rect 140759 457377 140827 457796
rect 127385 457211 134893 457333
rect 136832 457317 140827 457377
rect 127385 457049 127507 457211
rect 10720 456927 127507 457049
rect 134771 456973 134893 457211
rect 128832 456791 132834 456858
rect 134771 456851 142279 456973
rect 128832 456434 128913 456791
rect 10238 456233 128913 456434
rect 132752 456233 132834 456791
rect 10238 456148 132834 456233
rect 5343 455031 6129 455115
rect 8982 448336 133414 448422
rect 8982 446702 9147 448336
rect 10216 448269 133414 448336
rect 10216 446760 129000 448269
rect 132676 446760 133414 448269
rect 10216 446702 133414 446760
rect 8982 446610 133414 446702
rect 6463 439503 6744 439504
rect 6462 439485 6744 439503
rect 6462 438897 6476 439485
rect 6728 438897 6744 439485
rect 6462 438880 6744 438897
rect 6463 437005 6744 438880
rect 7368 439002 7592 439029
rect 7368 438204 7391 439002
rect 7570 438204 7592 439002
rect 7368 438178 7592 438204
rect 6447 436988 6755 437005
rect 6447 436151 6459 436988
rect 6743 436151 6755 436988
rect 6447 436136 6755 436151
rect 2398 435733 4680 435889
rect 2398 435716 2427 435733
rect 1703 435690 2427 435716
rect 7418 434511 7549 438178
rect 13208 437642 14598 437666
rect 13208 437442 13238 437642
rect 14564 437442 14598 437642
rect 13208 437416 14598 437442
rect 13394 436761 14363 437416
rect 13382 436724 14416 436761
rect 13382 434895 13424 436724
rect 14366 434895 14416 436724
rect 13382 434848 14416 434895
rect 7418 434380 141773 434511
rect 136831 434133 140827 434200
rect 136831 433676 136929 434133
rect 10249 433457 136929 433676
rect 140750 433676 140827 434133
rect 140750 433457 140833 433676
rect 10249 433366 140833 433457
rect 10219 433124 141383 433246
rect 10226 432924 132846 432928
rect 10226 432842 132847 432924
rect 10226 432642 128909 432842
rect 128832 432251 128909 432642
rect 132750 432251 132847 432842
rect 128832 432179 132847 432251
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 6302 429814 7162 429877
rect 11637 428240 13660 428297
rect 11637 428190 11697 428240
rect 11379 427828 11697 428190
rect 13585 428190 13660 428240
rect 13585 427828 13661 428190
rect 11379 427786 13661 427828
rect 11637 427782 13660 427786
rect 4524 426575 4680 426577
rect 4484 426541 4759 426575
rect 4484 425868 4522 426541
rect 4717 425868 4759 426541
rect 4484 425830 4759 425868
rect 8087 384757 9234 384793
rect 8087 384475 8126 384757
rect 9182 384475 9234 384757
rect 8087 384441 9234 384475
rect 8490 383290 9178 383354
rect 8490 382858 8553 383290
rect 9115 382858 9178 383290
rect 1694 382780 2576 382812
rect 8490 382807 9178 382858
rect 1694 382608 1730 382780
rect 2548 382608 2576 382780
rect 1694 382578 2576 382608
rect 8167 382289 9436 382347
rect 8167 381897 8241 382289
rect 9368 381897 9436 382289
rect 8167 381846 9436 381897
rect 7571 379992 9262 380019
rect 7571 379740 7617 379992
rect 9223 379740 9262 379992
rect 7571 379709 9262 379740
rect 7070 379384 136285 379463
rect 6839 379263 8545 379268
rect 6839 379239 9272 379263
rect 6839 378984 7609 379239
rect 9228 378984 9272 379239
rect 6839 378960 9272 378984
rect 7566 378955 9272 378960
rect 13425 360329 135815 360419
rect 13425 350850 13515 360329
rect 13711 359987 135473 360077
rect 13711 351650 13801 359987
rect 14063 359639 135125 359729
rect 14063 352450 14153 359639
rect 62370 359282 134778 359382
rect 59776 359034 60384 359062
rect 59776 358268 59802 359034
rect 60356 358268 60384 359034
rect 59776 358236 60384 358268
rect 62370 357580 62470 359282
rect 61740 357480 62470 357580
rect 62658 358928 134424 359028
rect 62658 356580 62758 358928
rect 61612 356480 62758 356580
rect 63062 358592 134088 358692
rect 63062 355580 63162 358592
rect 61612 355480 63162 355580
rect 63382 358220 133716 358320
rect 63382 354580 63482 358220
rect 61636 354480 63482 354580
rect 63680 357796 133292 357896
rect 63680 353580 63780 357796
rect 61702 353480 63780 353580
rect 63946 357476 132972 357576
rect 63946 352580 64046 357476
rect 61736 352480 64046 352580
rect 14063 352360 15233 352450
rect 13711 351560 15211 351650
rect 13425 350760 15111 350850
rect 4957 344582 5920 344626
rect 4957 344467 4993 344582
rect 5879 344467 5920 344582
rect 4957 344428 5920 344467
rect 4935 339653 6035 339688
rect 1528 339574 2590 339613
rect 1528 339376 1564 339574
rect 2527 339376 2590 339574
rect 1528 339348 2590 339376
rect 4935 339220 4983 339653
rect 5982 339220 6035 339653
rect 4935 339168 6035 339220
rect 2937 327203 3264 335928
rect 7718 335437 8004 336324
rect 8442 336159 9430 336225
rect 6704 335356 8008 335437
rect 6704 334800 6789 335356
rect 7923 334800 8008 335356
rect 6704 334714 8008 334800
rect 4943 334449 5832 334464
rect 4943 334263 4974 334449
rect 5809 334263 5832 334449
rect 4943 334244 5832 334263
rect 2937 326876 3601 327203
rect 3274 314651 3601 326876
rect 3032 314581 3801 314651
rect 3032 311780 3091 314581
rect 3736 311780 3801 314581
rect 3032 311699 3801 311780
rect 3274 298709 3601 311699
rect 8208 302233 8310 335770
rect 8442 335696 8496 336159
rect 9359 335696 9430 336159
rect 8442 335630 9430 335696
rect 11825 302878 12095 302887
rect 11825 302864 11839 302878
rect 10985 302801 11839 302864
rect 8208 302131 10338 302233
rect 5372 301415 6335 301432
rect 5372 301251 5395 301415
rect 6315 301251 6335 301415
rect 5372 301234 6335 301251
rect 5194 296534 6467 296612
rect 1917 296389 2979 296430
rect 1917 296191 1959 296389
rect 2922 296191 2979 296389
rect 1917 296165 2979 296191
rect 5194 296044 5290 296534
rect 6335 296044 6467 296534
rect 5194 295966 6467 296044
rect 8863 293051 9807 293093
rect 7037 292119 8427 292167
rect 7037 291597 7102 292119
rect 8352 291597 8427 292119
rect 7037 291557 8427 291597
rect 5372 291271 6070 291289
rect 5372 291105 5396 291271
rect 6049 291105 6070 291271
rect 5372 291088 6070 291105
rect 8647 290719 8716 292519
rect 8863 292471 8908 293051
rect 9750 292471 9807 293051
rect 8863 292434 9807 292471
rect 8647 290650 10169 290719
rect 8738 215318 8797 284463
rect 10100 215680 10169 290650
rect 10269 215849 10338 302131
rect 10985 285560 11048 302801
rect 11825 302797 11839 302801
rect 12083 302797 12095 302878
rect 11825 302787 12095 302797
rect 11825 302677 12092 302686
rect 11825 302671 11835 302677
rect 11153 302608 11835 302671
rect 11153 286561 11216 302608
rect 11825 302596 11835 302608
rect 12079 302596 12092 302677
rect 11825 302587 12092 302596
rect 11135 286547 11237 286561
rect 11135 286351 11151 286547
rect 11227 286351 11237 286547
rect 11135 286333 11237 286351
rect 10965 285546 11073 285560
rect 10965 285344 10980 285546
rect 11060 285344 11073 285546
rect 10965 285328 11073 285344
rect 10985 285319 11048 285328
rect 10269 215780 126517 215849
rect 10100 215611 126348 215680
rect 8738 215259 126044 215318
rect 8977 85362 9957 91084
rect 10673 89075 11473 89153
rect 10673 88436 10745 89075
rect 11391 88436 11473 89075
rect 10673 88355 11473 88436
rect 12383 89075 13183 89153
rect 12383 88436 12471 89075
rect 13117 88436 13183 89075
rect 12383 88355 13183 88436
rect 11007 85908 11127 88355
rect 12711 86343 12831 88355
rect 13018 88353 13183 88355
rect 12711 86223 125837 86343
rect 11007 85788 125468 85908
rect 8977 84367 9045 85362
rect 9901 84367 9957 85362
rect 8977 84275 9957 84367
rect 3503 44764 4633 44867
rect 3503 44203 3580 44764
rect 4529 44203 4633 44764
rect 3503 44125 4633 44203
rect 5595 44369 5844 44392
rect 3511 43657 3915 44125
rect 5595 44084 5614 44369
rect 5821 44143 5844 44369
rect 5821 44084 18729 44143
rect 5595 44063 18729 44084
rect 1456 39496 1714 39528
rect 1456 38894 1484 39496
rect 1684 38894 1714 39496
rect 1456 38866 1714 38894
rect 5652 39422 6511 39493
rect 5652 38923 5712 39422
rect 6434 38923 6511 39422
rect 18649 39010 18729 44063
rect 76611 39010 76691 42357
rect 18646 38930 76691 39010
rect 5652 38883 6511 38923
rect 76611 38916 76691 38930
rect 9094 35996 9417 36046
rect 8367 33414 8653 35650
rect 8853 34283 8923 35511
rect 9094 35396 9153 35996
rect 9363 35396 9417 35996
rect 17380 35877 34661 35893
rect 17380 35823 123139 35877
rect 9094 35350 9417 35396
rect 17394 34283 17464 35823
rect 34591 35807 123139 35823
rect 8853 34213 17464 34283
rect 60375 34705 60456 34715
rect 60375 34422 60381 34705
rect 60444 34422 60456 34705
rect 9065 33908 9908 33954
rect 9065 33660 9132 33908
rect 9845 33660 9908 33908
rect 9065 33610 9908 33660
rect 8220 33376 8803 33414
rect 8220 33163 8266 33376
rect 8753 33163 8803 33376
rect 8220 33133 8803 33163
rect 8367 33124 8653 33133
rect 9077 32717 9878 33610
rect 9069 32667 9912 32717
rect 9069 32419 9136 32667
rect 9849 32419 9912 32667
rect 9069 32373 9912 32419
rect 7204 28409 7656 28442
rect 7204 27214 7258 28409
rect 7592 27214 7656 28409
rect 60375 27699 60456 34422
rect 60535 34705 60616 34715
rect 60535 34422 60541 34705
rect 60604 34422 60616 34705
rect 60535 27859 60616 34422
rect 60695 34705 60776 34715
rect 60695 34422 60701 34705
rect 60764 34422 60776 34705
rect 60695 28019 60776 34422
rect 60855 34705 60936 34715
rect 60855 34422 60861 34705
rect 60924 34422 60936 34705
rect 60855 28179 60936 34422
rect 61015 34705 61096 34715
rect 61015 34422 61021 34705
rect 61084 34422 61096 34705
rect 61015 28339 61096 34422
rect 61175 34705 61256 34715
rect 61175 34422 61181 34705
rect 61244 34422 61256 34705
rect 61175 28499 61256 34422
rect 61335 34705 61416 34715
rect 61335 34422 61341 34705
rect 61404 34422 61416 34705
rect 61335 28659 61416 34422
rect 61495 34705 61576 34715
rect 61495 34422 61501 34705
rect 61564 34422 61576 34705
rect 61495 28819 61576 34422
rect 65251 34661 65332 34672
rect 65251 34421 65259 34661
rect 65322 34421 65332 34661
rect 65251 29471 65332 34421
rect 65411 34661 65492 34672
rect 65411 34421 65419 34661
rect 65482 34421 65492 34661
rect 65411 29631 65492 34421
rect 65571 34661 65652 34672
rect 65571 34421 65579 34661
rect 65642 34421 65652 34661
rect 65571 29791 65652 34421
rect 65731 34661 65812 34672
rect 65731 34421 65739 34661
rect 65802 34421 65812 34661
rect 65731 29951 65812 34421
rect 65891 34661 65972 34672
rect 65891 34421 65899 34661
rect 65962 34421 65972 34661
rect 65891 30111 65972 34421
rect 66051 34661 66132 34672
rect 66051 34421 66059 34661
rect 66122 34421 66132 34661
rect 66051 30271 66132 34421
rect 66211 34661 66292 34672
rect 66211 34421 66219 34661
rect 66282 34421 66292 34661
rect 66211 30431 66292 34421
rect 66371 34661 66452 34672
rect 66371 34421 66379 34661
rect 66442 34421 66452 34661
rect 66371 30591 66452 34421
rect 66371 30510 120519 30591
rect 66211 30350 120359 30431
rect 66051 30190 120199 30271
rect 65891 30030 120039 30111
rect 65731 29870 119879 29951
rect 65571 29710 119719 29791
rect 65411 29550 119559 29631
rect 65251 29390 119399 29471
rect 61495 28738 118747 28819
rect 61335 28578 118587 28659
rect 61175 28418 118427 28499
rect 61015 28258 118267 28339
rect 60855 28098 118107 28179
rect 60695 27938 117947 28019
rect 60535 27778 117787 27859
rect 60375 27618 117627 27699
rect 7204 27149 7656 27214
rect 117546 3735 117627 27618
rect 117706 3895 117787 27778
rect 117866 4055 117947 27938
rect 118026 4215 118107 28098
rect 118186 4375 118267 28258
rect 118346 4535 118427 28418
rect 118506 4695 118587 28578
rect 118666 4855 118747 28738
rect 119318 5507 119399 29390
rect 119478 5667 119559 29550
rect 119638 5827 119719 29710
rect 119798 5987 119879 29870
rect 119958 6147 120039 30030
rect 120118 6307 120199 30190
rect 120278 6467 120359 30350
rect 120438 6627 120519 30510
rect 123069 7693 123139 35807
rect 125348 8065 125468 85788
rect 125717 8469 125837 86223
rect 125985 8631 126044 215259
rect 126279 8829 126348 215611
rect 126448 8998 126517 215780
rect 132872 11398 132972 357476
rect 133192 11794 133292 357796
rect 133616 12132 133716 358220
rect 133988 12472 134088 358592
rect 134324 12866 134424 358928
rect 134678 13348 134778 359282
rect 135035 13783 135125 359639
rect 135383 14233 135473 359987
rect 135725 14607 135815 360329
rect 136206 14933 136285 379384
rect 141261 15423 141383 433124
rect 141642 15813 141773 434380
rect 142157 16319 142279 456851
rect 142468 16608 142568 476633
rect 263426 476584 263662 477313
rect 265591 476584 265741 477313
rect 263426 476391 265741 476584
rect 245574 473106 247889 473256
rect 245574 472377 245788 473106
rect 247717 472377 247889 473106
rect 245574 472184 247889 472377
rect 279035 463726 282207 463786
rect 263426 384713 265741 384863
rect 263426 383984 263662 384713
rect 265591 383984 265741 384713
rect 263426 383791 265741 383984
rect 245574 383106 247889 383256
rect 245574 382377 245788 383106
rect 247717 382377 247889 383106
rect 245574 382184 247889 382377
rect 279035 373726 281927 373786
rect 263426 294713 265741 294863
rect 263426 293984 263662 294713
rect 265591 293984 265741 294713
rect 263426 293791 265741 293984
rect 245574 293106 247889 293256
rect 245574 292377 245788 293106
rect 247717 292377 247889 293106
rect 245574 292184 247889 292377
rect 279035 283726 281647 283786
rect 263426 204713 265741 204863
rect 263426 203984 263662 204713
rect 265591 203984 265741 204713
rect 263426 203791 265741 203984
rect 245574 203106 247889 203256
rect 245574 202377 245788 203106
rect 247717 202377 247889 203106
rect 245574 202184 247889 202377
rect 279035 193726 281367 193786
rect 263426 114713 265741 114863
rect 263426 113984 263662 114713
rect 265591 113984 265741 114713
rect 263426 113791 265741 113984
rect 245574 113106 247889 113256
rect 245574 112377 245788 113106
rect 247717 112377 247889 113106
rect 245574 112184 247889 112377
rect 279035 103726 281087 103786
rect 142468 16508 257918 16608
rect 142157 16197 254401 16319
rect 141642 15682 250832 15813
rect 141261 15301 247289 15423
rect 181943 14965 182423 14982
rect 181943 14933 181967 14965
rect 136206 14869 181967 14933
rect 182409 14869 182423 14965
rect 136206 14855 182423 14869
rect 136206 14854 182413 14855
rect 135725 14517 243735 14607
rect 135383 14143 240199 14233
rect 135035 13693 236651 13783
rect 134678 13248 233096 13348
rect 134324 12766 229548 12866
rect 133988 12372 226022 12472
rect 133616 12032 222474 12132
rect 133192 11694 218936 11794
rect 132872 11298 215378 11398
rect 126448 8929 208280 8998
rect 126279 8760 204722 8829
rect 125985 8572 201171 8631
rect 125717 8379 197644 8469
rect 125348 7975 194083 8065
rect 123069 7623 190531 7693
rect 181525 7436 182295 7460
rect 181525 7340 181554 7436
rect 182266 7423 182295 7436
rect 182266 7342 187002 7423
rect 182266 7340 182295 7342
rect 181525 7316 182295 7340
rect 120438 6546 183462 6627
rect 120278 6386 179898 6467
rect 120118 6226 176347 6307
rect 119958 6066 172808 6147
rect 119798 5906 169281 5987
rect 119638 5746 165717 5827
rect 119478 5586 162172 5667
rect 119318 5426 158633 5507
rect 118666 4774 155075 4855
rect 118506 4614 151523 4695
rect 118346 4454 147997 4535
rect 118186 4294 144439 4375
rect 118026 4134 140906 4215
rect 117866 3974 137348 4055
rect 117706 3814 133803 3895
rect 117546 3654 130270 3735
rect 130189 1280 130270 3654
rect 133722 1280 133803 3814
rect 137267 1280 137348 3974
rect 140825 1280 140906 4134
rect 144358 1280 144439 4294
rect 147916 1280 147997 4454
rect 151442 1280 151523 4614
rect 154994 1280 155075 4774
rect 158552 1280 158633 5426
rect 162091 1280 162172 5586
rect 165636 1280 165717 5746
rect 169200 1296 169281 5906
rect 169200 1280 169280 1296
rect 172727 1280 172808 6066
rect 176266 1280 176347 6226
rect 179817 1280 179898 6386
rect 183381 1280 183462 6546
rect 186921 1280 187002 7342
rect 190461 1280 190531 7623
rect 193993 1280 194083 7975
rect 197554 1280 197644 8379
rect 201112 1280 201171 8572
rect 204653 1280 204722 8760
rect 208211 1280 208280 8929
rect 215278 1280 215378 11298
rect 218836 1296 218936 11694
rect 222374 1296 222474 12032
rect 225922 1296 226022 12372
rect 218836 1280 218924 1296
rect 222374 1280 222470 1296
rect 225922 1280 226016 1296
rect 229448 1280 229548 12766
rect 232996 1280 233096 13248
rect 236561 1280 236651 13693
rect 240109 1280 240199 14143
rect 243645 1280 243735 14517
rect 247167 1280 247289 15301
rect 250701 1280 250832 15682
rect 254279 1296 254401 16197
rect 254279 1280 254384 1296
rect 257818 1280 257918 16508
rect 261092 9685 261152 11294
rect 264640 9812 264700 11294
rect 268188 9942 268248 11294
rect 271736 10070 271796 11294
rect 275284 10196 275344 11294
rect 278214 10324 278274 11294
rect 278562 10452 278622 11294
rect 278910 10582 278970 11294
rect 279258 10709 279318 11294
rect 279606 10837 279666 11294
rect 279954 10965 280014 11294
rect 280302 11093 280362 11294
rect 280227 11088 280448 11093
rect 280227 11032 280236 11088
rect 280439 11032 280448 11088
rect 280227 11027 280448 11032
rect 279879 10960 280100 10965
rect 279879 10904 279888 10960
rect 280091 10904 280100 10960
rect 279879 10899 280100 10904
rect 279510 10832 279731 10837
rect 279510 10776 279573 10832
rect 279722 10776 279731 10832
rect 279510 10771 279731 10776
rect 279186 10704 279407 10709
rect 279186 10648 279262 10704
rect 279398 10648 279407 10704
rect 279186 10643 279407 10648
rect 278837 10577 279058 10582
rect 278837 10521 278859 10577
rect 279049 10521 279058 10577
rect 278837 10516 279058 10521
rect 278479 10447 278700 10452
rect 278479 10391 278570 10447
rect 278691 10391 278700 10447
rect 278479 10386 278700 10391
rect 278145 10319 278366 10324
rect 278145 10263 278154 10319
rect 278357 10263 278366 10319
rect 278145 10258 278366 10263
rect 275208 10191 275429 10196
rect 275208 10135 275217 10191
rect 275420 10135 275429 10191
rect 275208 10130 275429 10135
rect 271654 10065 271878 10070
rect 271654 10009 271663 10065
rect 271866 10009 271878 10065
rect 271654 10004 271878 10009
rect 268130 9937 268351 9942
rect 268130 9881 268139 9937
rect 268342 9881 268351 9937
rect 268130 9876 268351 9881
rect 264553 9807 264774 9812
rect 264553 9751 264562 9807
rect 264765 9751 264774 9807
rect 264553 9746 264774 9751
rect 261008 9680 261229 9685
rect 261008 9624 261017 9680
rect 261220 9624 261229 9680
rect 261008 9619 261229 9624
rect 261092 7841 261152 9619
rect 264640 8091 264700 9746
rect 268188 8330 268248 9876
rect 271736 8569 271796 10004
rect 275284 8842 275344 10130
rect 275284 8782 275627 8842
rect 271736 8509 272079 8569
rect 268188 8270 268532 8330
rect 264640 8031 264996 8091
rect 261092 7781 261448 7841
rect 261388 1280 261448 7781
rect 264936 1280 264996 8031
rect 268472 1280 268532 8270
rect 272019 1280 272079 8509
rect 275567 1280 275627 8782
rect 278214 3103 278274 10258
rect 278562 3410 278622 10386
rect 278910 3660 278970 10516
rect 279258 3967 279318 10643
rect 279606 4320 279666 10771
rect 279954 4581 280014 10899
rect 280302 4820 280362 11027
rect 281027 5033 281087 103726
rect 281307 5313 281367 193726
rect 281587 5593 281647 283726
rect 281867 5873 281927 373726
rect 282147 6153 282207 463726
rect 282427 6433 282487 553726
rect 282707 6713 282767 643726
rect 303962 643726 307687 643786
rect 286531 281299 286590 281335
rect 286531 9685 286590 281121
rect 298623 281284 298693 281337
rect 286731 280629 286790 280703
rect 286731 9813 286790 280434
rect 286931 279501 286990 279594
rect 286931 9941 286990 279306
rect 287131 277413 287190 277500
rect 287131 10069 287190 277218
rect 287331 275318 287390 275460
rect 287331 10198 287390 275123
rect 287531 273227 287590 273300
rect 287531 10325 287590 273032
rect 287731 270055 287790 270136
rect 287731 10453 287790 269860
rect 287931 264802 287990 264864
rect 287931 10581 287990 264595
rect 298423 264296 298493 264355
rect 298223 208190 298293 208297
rect 288131 197629 288190 197695
rect 288131 10709 288190 197431
rect 298023 155592 298093 155657
rect 297823 103096 297893 103167
rect 288309 87253 288390 87280
rect 288309 87009 288390 87051
rect 288331 10837 288390 87009
rect 288552 79955 288870 80019
rect 288552 10965 288616 79955
rect 297459 68899 297693 68969
rect 288910 47431 289456 47493
rect 288910 11093 288972 47431
rect 297246 46310 297494 46449
rect 290073 30905 290992 30949
rect 290073 30361 290122 30905
rect 290933 30361 290992 30905
rect 290073 30317 290992 30361
rect 288826 11088 289047 11093
rect 288826 11032 288835 11088
rect 289038 11032 289047 11088
rect 288826 11027 289047 11032
rect 288452 10960 288673 10965
rect 288452 10904 288461 10960
rect 288664 10904 288673 10960
rect 288452 10899 288673 10904
rect 288248 10832 288469 10837
rect 288248 10776 288257 10832
rect 288460 10776 288469 10832
rect 288248 10771 288469 10776
rect 288053 10704 288274 10709
rect 288053 10648 288062 10704
rect 288265 10648 288274 10704
rect 288053 10643 288274 10648
rect 287856 10576 288077 10581
rect 287856 10520 287865 10576
rect 288068 10520 288077 10576
rect 287856 10515 288077 10520
rect 287654 10448 287875 10453
rect 287654 10392 287663 10448
rect 287866 10392 287875 10448
rect 287654 10387 287875 10392
rect 287455 10320 287676 10325
rect 287455 10264 287464 10320
rect 287667 10264 287676 10320
rect 287455 10259 287676 10264
rect 287246 10193 287467 10198
rect 287246 10137 287255 10193
rect 287458 10137 287467 10193
rect 287246 10132 287467 10137
rect 287060 10064 287281 10069
rect 287060 10008 287069 10064
rect 287272 10008 287281 10064
rect 287060 10003 287281 10008
rect 286857 9936 287078 9941
rect 286857 9880 286866 9936
rect 287069 9880 287078 9936
rect 286857 9875 287078 9880
rect 286670 9808 286891 9813
rect 286670 9752 286679 9808
rect 286882 9752 286891 9808
rect 286670 9747 286891 9752
rect 286452 9680 286673 9685
rect 286452 9624 286461 9680
rect 286664 9624 286673 9680
rect 286452 9619 286673 9624
rect 286531 9520 286590 9619
rect 286731 9520 286790 9747
rect 286931 9520 286990 9875
rect 287131 9520 287190 10003
rect 287331 9520 287390 10132
rect 287531 9520 287590 10259
rect 287731 9520 287790 10387
rect 287931 9520 287990 10515
rect 288131 9520 288190 10643
rect 288331 9520 288390 10771
rect 288552 9520 288616 10899
rect 288910 9520 288972 11027
rect 297423 10535 297493 46310
rect 297350 10530 297571 10535
rect 297350 10474 297359 10530
rect 297562 10474 297571 10530
rect 297350 10469 297571 10474
rect 297423 9617 297493 10469
rect 297623 10407 297693 68899
rect 297546 10402 297767 10407
rect 297546 10346 297555 10402
rect 297758 10346 297767 10402
rect 297546 10341 297767 10346
rect 297623 9617 297693 10341
rect 297823 10279 297893 102891
rect 297744 10274 297965 10279
rect 297744 10218 297753 10274
rect 297956 10218 297965 10274
rect 297744 10213 297965 10218
rect 297823 9617 297893 10213
rect 298023 10150 298093 155388
rect 297951 10145 298172 10150
rect 297951 10089 297960 10145
rect 298163 10089 298172 10145
rect 297951 10084 298172 10089
rect 298023 9617 298093 10084
rect 298223 10023 298293 207988
rect 298149 10018 298370 10023
rect 298149 9962 298158 10018
rect 298361 9962 298370 10018
rect 298149 9957 298370 9962
rect 298223 9617 298293 9957
rect 298423 9895 298493 264095
rect 298345 9890 298566 9895
rect 298345 9834 298354 9890
rect 298557 9834 298566 9890
rect 298345 9829 298566 9834
rect 298423 9617 298493 9829
rect 298623 9767 298693 281046
rect 298862 57142 298998 57176
rect 298862 56610 298894 57142
rect 298962 56610 298998 57142
rect 298862 56584 298998 56610
rect 298886 10694 298958 56584
rect 298868 10678 299194 10694
rect 298868 10620 298896 10678
rect 299168 10620 299194 10678
rect 298868 10600 299194 10620
rect 298886 10546 298958 10600
rect 298541 9762 298762 9767
rect 298541 9706 298550 9762
rect 298753 9706 298762 9762
rect 298541 9701 298762 9706
rect 298623 9617 298693 9701
rect 303962 7352 304022 643726
rect 444175 617823 448174 617824
rect 444175 617699 560181 617823
rect 444175 614087 444372 617699
rect 448011 614087 560181 617699
rect 444175 613931 560181 614087
rect 444223 613929 560181 613931
rect 513415 609778 520733 610315
rect 508780 594670 510602 595116
rect 513415 595070 513911 609778
rect 513414 594741 513911 595070
rect 513415 593259 513911 594741
rect 520276 593259 520733 609778
rect 556287 602040 560181 613929
rect 556287 601770 560183 602040
rect 556287 593934 556508 601770
rect 560007 595003 560183 601770
rect 560007 594682 569275 595003
rect 560007 593934 560183 594682
rect 556287 593698 560183 593934
rect 513415 592789 520733 593259
rect 568954 589367 569275 594682
rect 583563 589372 583751 589414
rect 568861 589315 569347 589367
rect 568861 588943 568944 589315
rect 569285 588943 569347 589315
rect 568861 588870 569347 588943
rect 583563 588859 583568 589372
rect 583746 588859 583751 589372
rect 583563 588791 583751 588859
rect 583568 587366 583746 588791
rect 563565 587188 583746 587366
rect 573463 586727 574467 586813
rect 573463 585613 573573 586727
rect 574366 585613 574467 586727
rect 573463 585534 574467 585613
rect 583830 584564 584262 584602
rect 583830 584260 583874 584564
rect 584212 584260 584262 584564
rect 583830 584232 584262 584260
rect 577087 584173 577726 584230
rect 577087 583409 577145 584173
rect 577661 583409 577726 584173
rect 577087 583360 577726 583409
rect 563548 582534 565009 582654
rect 510422 576926 518844 577547
rect 510422 570179 510907 576926
rect 518330 570179 518844 576926
rect 510422 569612 518844 570179
rect 556374 572886 560268 573078
rect 556374 566873 556611 572886
rect 452076 566724 556611 566873
rect 321050 564704 323365 564854
rect 321050 563975 321200 564704
rect 323129 563975 323365 564704
rect 321050 563782 323365 563975
rect 338902 563097 341217 563247
rect 338902 562368 339074 563097
rect 341003 562368 341217 563097
rect 452076 563112 452351 566724
rect 455990 563187 556611 566724
rect 560065 566873 560268 572886
rect 560065 565322 560278 566873
rect 560065 565066 562890 565322
rect 560065 564711 560571 565066
rect 562698 564711 562890 565066
rect 560065 564413 562890 564711
rect 560065 563187 560278 564413
rect 455990 563112 560278 563187
rect 452076 562979 560278 563112
rect 338902 562175 341217 562368
rect 438929 561647 439466 561660
rect 438929 561526 438947 561647
rect 439446 561643 439466 561647
rect 564895 561643 565009 582534
rect 565411 581852 565859 581897
rect 565411 581487 565447 581852
rect 565813 581758 565859 581852
rect 565813 581725 579385 581758
rect 565813 581498 578165 581725
rect 579312 581498 579385 581725
rect 565813 581487 579385 581498
rect 565411 581473 579385 581487
rect 565411 581449 565859 581473
rect 439446 561529 565009 561643
rect 566678 581140 579582 581228
rect 439446 561526 439466 561529
rect 438929 561509 439466 561526
rect 439337 561071 439874 561084
rect 439337 560950 439355 561071
rect 439854 561067 439874 561071
rect 439854 561044 439888 561067
rect 566678 561044 566766 581140
rect 568880 580907 579894 581000
rect 568880 580660 568964 580907
rect 567629 580543 567862 580597
rect 567629 579827 567667 580543
rect 567829 579827 567862 580543
rect 568892 580566 568964 580660
rect 569295 580660 579894 580907
rect 569295 580566 569368 580660
rect 568892 580524 569368 580566
rect 567629 579773 567862 579827
rect 439854 560956 566766 561044
rect 439854 560953 439888 560956
rect 439854 560950 439874 560953
rect 439337 560933 439874 560950
rect 422745 558959 423751 558994
rect 422745 558790 422782 558959
rect 423705 558926 423751 558959
rect 567690 558926 567807 579773
rect 423705 558809 567807 558926
rect 423705 558790 423751 558809
rect 422745 558762 423751 558790
rect 304242 553726 307687 553786
rect 304242 7746 304302 553726
rect 575990 498421 576687 498523
rect 575990 496743 576075 498421
rect 576616 496743 576687 498421
rect 575990 496650 576687 496743
rect 574914 496291 575907 496393
rect 574914 495447 575013 496291
rect 575808 495447 575907 496291
rect 574914 495358 575907 495447
rect 583438 495102 584234 495148
rect 576700 494849 577862 494922
rect 576700 493993 576790 494849
rect 577757 493993 577862 494849
rect 583438 494882 583490 495102
rect 584168 494882 584234 495102
rect 583438 494838 584234 494882
rect 576700 493929 577862 493993
rect 578266 492276 579461 492320
rect 578266 492070 578317 492276
rect 579412 492070 579461 492276
rect 578266 492032 579461 492070
rect 460166 491840 460662 491858
rect 460166 491736 460200 491840
rect 460638 491810 460662 491840
rect 460638 491736 579262 491810
rect 460166 491730 579262 491736
rect 460166 491710 460662 491730
rect 578225 491568 579451 491594
rect 578225 491321 578266 491568
rect 579420 491321 579451 491568
rect 578225 491282 579451 491321
rect 321050 474704 323365 474854
rect 321050 473975 321200 474704
rect 323129 473975 323365 474704
rect 321050 473782 323365 473975
rect 338902 473097 341217 473247
rect 338902 472368 339074 473097
rect 341003 472368 341217 473097
rect 338902 472175 341217 472368
rect 304522 463726 307687 463786
rect 304522 8078 304582 463726
rect 557755 435818 557986 435844
rect 557755 434769 557782 435818
rect 557961 434975 557986 435818
rect 557961 434769 559425 434975
rect 557755 434744 559425 434769
rect 582171 433815 583321 434170
rect 583433 433815 583444 434170
rect 582185 431416 583313 431771
rect 583425 431416 583453 431771
rect 419480 422228 421176 422253
rect 419480 422017 419509 422228
rect 421145 422188 421176 422228
rect 421145 422035 559381 422188
rect 421145 422017 421176 422035
rect 419480 421993 421176 422017
rect 452250 421269 559235 421330
rect 452250 421117 452329 421269
rect 452172 420738 452329 421117
rect 452250 420650 452329 420738
rect 456074 421117 559235 421269
rect 456074 420738 559442 421117
rect 456074 420650 559235 420738
rect 452250 420572 559235 420650
rect 444312 419339 559230 419413
rect 444312 419211 444386 419339
rect 444073 418832 444386 419211
rect 444312 418708 444386 418832
rect 447969 419211 559230 419339
rect 447969 418832 559373 419211
rect 447969 418708 559230 418832
rect 444312 418647 559230 418708
rect 553923 415365 554697 415400
rect 553923 415328 554002 415365
rect 456842 415208 554002 415328
rect 321050 384704 323365 384854
rect 321050 383975 321200 384704
rect 323129 383975 323365 384704
rect 321050 383782 323365 383975
rect 338902 383097 341217 383247
rect 338902 382368 339074 383097
rect 341003 382368 341217 383097
rect 338902 382175 341217 382368
rect 304802 373726 307687 373786
rect 304802 8398 304862 373726
rect 338902 295097 341217 295247
rect 338902 294368 339074 295097
rect 341003 294368 341217 295097
rect 338902 294175 341217 294368
rect 321062 292916 323377 293065
rect 321062 292187 321212 292916
rect 323141 292187 323377 292916
rect 321062 291994 323377 292187
rect 305082 283726 307687 283786
rect 305082 8711 305142 283726
rect 439358 216572 439534 216600
rect 439358 216140 439388 216572
rect 439512 216270 439534 216572
rect 439512 216150 456536 216270
rect 439512 216140 439534 216150
rect 439358 216120 439534 216140
rect 321050 204704 323365 204854
rect 321050 203975 321200 204704
rect 323129 203975 323365 204704
rect 321050 203782 323365 203975
rect 338902 203097 341217 203247
rect 338902 202368 339074 203097
rect 341003 202368 341217 203097
rect 338902 202175 341217 202368
rect 305362 193726 307687 193786
rect 305362 9043 305422 193726
rect 321050 114704 323365 114854
rect 321050 113975 321200 114704
rect 323129 113975 323365 114704
rect 321050 113782 323365 113975
rect 338902 113097 341217 113247
rect 338902 112368 339074 113097
rect 341003 112368 341217 113097
rect 338902 112175 341217 112368
rect 305642 103726 307687 103786
rect 305642 9401 305702 103726
rect 456416 15774 456536 216150
rect 456270 15732 456558 15774
rect 456270 14942 456314 15732
rect 456522 14942 456558 15732
rect 456270 14892 456558 14942
rect 403228 10535 403288 10593
rect 403147 10530 403368 10535
rect 403147 10474 403156 10530
rect 403359 10474 403368 10530
rect 403147 10469 403368 10474
rect 305642 9341 399747 9401
rect 305362 8983 392663 9043
rect 305082 8651 385566 8711
rect 304802 8338 378475 8398
rect 304522 8018 371358 8078
rect 304242 7686 364274 7746
rect 303962 7292 357200 7352
rect 282707 6653 346571 6713
rect 282427 6373 339462 6433
rect 282147 6093 332374 6153
rect 281867 5813 325275 5873
rect 281587 5533 318187 5593
rect 281307 5253 311088 5313
rect 281027 4973 304000 5033
rect 280302 4760 300447 4820
rect 279954 4521 296911 4581
rect 279606 4260 293364 4320
rect 279258 3907 289816 3967
rect 278910 3600 286269 3660
rect 278562 3350 282721 3410
rect 278214 3043 279174 3103
rect 279114 1280 279174 3043
rect 282661 1280 282721 3350
rect 286209 1280 286269 3600
rect 289756 1280 289816 3907
rect 293304 1280 293364 4260
rect 296851 1280 296911 4521
rect 300387 1280 300447 4760
rect 303940 1280 304000 4973
rect 311028 1280 311088 5253
rect 318127 1280 318187 5533
rect 325215 1280 325275 5813
rect 332314 1280 332374 6093
rect 339402 1280 339462 6373
rect 346511 1280 346571 6653
rect 357140 1280 357200 7292
rect 364214 1280 364274 7686
rect 371298 1280 371358 8018
rect 378415 1280 378475 8338
rect 385506 1280 385566 8651
rect 392603 1280 392663 8983
rect 399687 1280 399747 9341
rect 403228 1280 403288 10469
rect 406776 10407 406836 10593
rect 406701 10402 406922 10407
rect 406701 10346 406710 10402
rect 406913 10346 406922 10402
rect 406701 10341 406922 10346
rect 406776 1280 406836 10341
rect 410324 10279 410384 10593
rect 410259 10274 410480 10279
rect 410259 10218 410268 10274
rect 410471 10218 410480 10274
rect 410259 10213 410480 10218
rect 410324 1280 410384 10213
rect 413872 10149 413932 10593
rect 413807 10144 414028 10149
rect 413807 10088 413816 10144
rect 414019 10088 414028 10144
rect 413807 10083 414028 10088
rect 413872 1280 413932 10083
rect 417420 10022 417480 10593
rect 417344 10017 417565 10022
rect 417344 9961 417353 10017
rect 417556 9961 417565 10017
rect 417344 9956 417565 9961
rect 417420 1280 417480 9956
rect 420968 9893 421028 10593
rect 420880 9888 421101 9893
rect 420880 9832 420889 9888
rect 421092 9832 421101 9888
rect 420880 9827 421101 9832
rect 420968 1280 421028 9827
rect 424516 9766 424576 10593
rect 424454 9761 424675 9766
rect 424454 9705 424463 9761
rect 424666 9705 424675 9761
rect 424454 9700 424675 9705
rect 424516 1280 424576 9700
rect 456842 7086 456962 415208
rect 553923 415181 554002 415208
rect 554622 415181 554697 415365
rect 553923 415145 554697 415181
rect 556073 415373 556847 415414
rect 556073 415189 556144 415373
rect 556764 415328 556847 415373
rect 556764 415208 559384 415328
rect 556764 415189 556847 415208
rect 556073 415159 556847 415189
rect 553923 414625 554697 414660
rect 428023 6966 456962 7086
rect 457161 414588 477255 414609
rect 553923 414588 554002 414625
rect 457161 414489 554002 414588
rect 428023 1296 428143 6966
rect 457161 6473 457281 414489
rect 477058 414468 554002 414489
rect 553923 414441 554002 414468
rect 554622 414441 554697 414625
rect 553923 414405 554697 414441
rect 556073 414633 556847 414674
rect 556073 414449 556144 414633
rect 556764 414588 556847 414633
rect 556764 414468 559484 414588
rect 556764 414449 556847 414468
rect 556073 414419 556847 414449
rect 547144 413369 559324 413371
rect 431556 6353 457281 6473
rect 458295 412900 458412 412928
rect 1324 800 1436 1280
rect 2506 800 2618 1280
rect 3688 800 3800 1280
rect 4870 800 4982 1280
rect 6052 800 6164 1280
rect 7234 800 7346 1280
rect 8416 800 8528 1280
rect 9598 800 9710 1280
rect 10780 800 10892 1280
rect 11962 800 12074 1280
rect 13144 800 13256 1280
rect 14326 800 14438 1280
rect 15508 800 15620 1280
rect 16690 800 16802 1280
rect 17872 800 17984 1280
rect 19054 800 19166 1280
rect 20236 800 20348 1280
rect 21418 800 21530 1280
rect 22600 800 22712 1280
rect 23782 800 23894 1280
rect 24964 800 25076 1280
rect 26146 800 26258 1280
rect 27328 800 27440 1280
rect 28510 800 28622 1280
rect 29692 800 29804 1280
rect 30874 800 30986 1280
rect 32056 800 32168 1280
rect 33238 800 33350 1280
rect 34420 800 34532 1280
rect 35602 800 35714 1280
rect 36784 800 36896 1280
rect 37966 800 38078 1280
rect 39148 800 39260 1280
rect 40330 800 40442 1280
rect 41512 800 41624 1280
rect 42694 800 42806 1280
rect 43876 800 43988 1280
rect 45058 800 45170 1280
rect 46240 800 46352 1280
rect 47422 800 47534 1280
rect 48604 800 48716 1280
rect 49786 800 49898 1280
rect 50968 800 51080 1280
rect 52150 800 52262 1280
rect 53332 800 53444 1280
rect 54514 800 54626 1280
rect 55696 800 55808 1280
rect 56878 800 56990 1280
rect 58060 800 58172 1280
rect 59242 800 59354 1280
rect 60424 800 60536 1280
rect 61606 800 61718 1280
rect 62788 800 62900 1280
rect 63970 800 64082 1280
rect 65152 800 65264 1280
rect 66334 800 66446 1280
rect 67516 800 67628 1280
rect 68698 800 68810 1280
rect 69880 800 69992 1280
rect 71062 800 71174 1280
rect 72244 800 72356 1280
rect 73426 800 73538 1280
rect 74608 800 74720 1280
rect 75790 800 75902 1280
rect 76972 800 77084 1280
rect 78154 800 78266 1280
rect 79336 800 79448 1280
rect 80518 800 80630 1280
rect 81700 800 81812 1280
rect 82882 800 82994 1280
rect 84064 800 84176 1280
rect 85246 800 85358 1280
rect 86428 800 86540 1280
rect 87610 800 87722 1280
rect 88792 800 88904 1280
rect 89974 800 90086 1280
rect 91156 800 91268 1280
rect 92338 800 92450 1280
rect 93520 800 93632 1280
rect 94702 800 94814 1280
rect 95884 800 95996 1280
rect 97066 800 97178 1280
rect 98248 800 98360 1280
rect 99430 800 99542 1280
rect 100612 800 100724 1280
rect 101794 800 101906 1280
rect 102976 800 103088 1280
rect 104158 800 104270 1280
rect 105340 800 105452 1280
rect 106522 800 106634 1280
rect 107704 800 107816 1280
rect 108886 800 108998 1280
rect 110068 800 110180 1279
rect 111250 800 111362 1280
rect 112432 800 112544 1280
rect 113614 800 113726 1280
rect 114796 800 114908 1280
rect 115978 800 116090 1280
rect 117160 800 117272 1280
rect 118342 800 118454 1280
rect 119524 800 119636 1280
rect 120706 800 120818 1280
rect 121888 800 122000 1280
rect 123070 800 123182 1280
rect 124252 800 124364 1280
rect 125434 800 125546 1280
rect 126616 0 126728 1280
rect 127798 0 127910 1280
rect 128980 800 129092 1280
rect 130162 0 130274 1280
rect 131344 0 131456 1280
rect 132526 800 132638 1280
rect 133708 0 133820 1280
rect 134890 0 135002 1280
rect 136072 800 136184 1280
rect 137254 0 137366 1280
rect 138436 0 138548 1280
rect 139618 800 139730 1279
rect 140800 0 140912 1280
rect 141982 0 142094 1280
rect 143164 800 143276 1279
rect 144346 0 144458 1280
rect 145528 1279 145640 1280
rect 145528 1178 145648 1279
rect 145528 0 145640 1178
rect 146710 800 146822 1279
rect 147892 0 148004 1280
rect 149074 0 149186 1280
rect 150256 800 150368 1279
rect 151438 0 151550 1280
rect 152620 0 152732 1280
rect 153802 800 153914 1279
rect 154984 0 155096 1280
rect 156166 0 156278 1280
rect 157348 800 157460 1279
rect 158530 0 158642 1280
rect 159712 1279 159824 1280
rect 159712 1152 159836 1279
rect 159712 0 159824 1152
rect 160894 800 161006 1279
rect 162076 0 162188 1280
rect 163258 1279 163370 1280
rect 163258 1108 163374 1279
rect 163258 0 163370 1108
rect 164440 800 164552 1279
rect 165622 0 165734 1280
rect 166804 1279 166916 1280
rect 166804 1140 166922 1279
rect 166804 0 166916 1140
rect 167986 800 168098 1279
rect 169168 0 169280 1280
rect 170350 1112 170464 1280
rect 170350 0 170462 1112
rect 171532 800 171644 1279
rect 172714 0 172826 1280
rect 173896 0 174008 1280
rect 175078 800 175190 1279
rect 176260 0 176372 1280
rect 177442 0 177554 1280
rect 178624 800 178736 1279
rect 179806 0 179918 1280
rect 180988 0 181100 1280
rect 182170 800 182282 1279
rect 183352 0 183464 1280
rect 184534 0 184646 1280
rect 185716 800 185828 1279
rect 186898 0 187010 1280
rect 188080 0 188192 1280
rect 189262 800 189374 1279
rect 190444 0 190556 1280
rect 191626 0 191738 1280
rect 192808 800 192920 1279
rect 193990 0 194102 1280
rect 195172 0 195284 1280
rect 196354 800 196466 1279
rect 197536 0 197648 1280
rect 198718 0 198830 1280
rect 199900 800 200012 1280
rect 201082 0 201194 1280
rect 202264 0 202376 1280
rect 203446 800 203558 1280
rect 204628 0 204740 1280
rect 205810 0 205922 1280
rect 206992 800 207104 1280
rect 208174 0 208286 1280
rect 209356 0 209468 1280
rect 210538 800 210650 1280
rect 211720 0 211832 1280
rect 212902 0 213014 1280
rect 214084 800 214196 1280
rect 215266 0 215378 1280
rect 217630 800 217742 1280
rect 218812 0 218924 1280
rect 219994 0 220106 1279
rect 221176 800 221288 1280
rect 222358 0 222470 1280
rect 223540 0 223652 1279
rect 224722 800 224834 1280
rect 225904 0 226016 1280
rect 227086 0 227198 1279
rect 228268 800 228380 1280
rect 229448 1279 229562 1280
rect 229450 0 229562 1279
rect 230632 0 230744 1280
rect 231814 800 231926 1280
rect 232996 0 233108 1280
rect 234178 0 234290 1280
rect 235360 800 235472 1280
rect 236542 0 236654 1280
rect 237724 0 237836 1280
rect 238906 800 239018 1280
rect 240088 0 240200 1280
rect 241270 0 241382 1280
rect 242452 800 242564 1280
rect 243634 0 243746 1280
rect 244816 0 244928 1280
rect 245998 800 246110 1280
rect 247180 0 247292 1280
rect 248362 0 248474 1280
rect 249544 800 249656 1280
rect 250726 0 250838 1280
rect 251908 0 252020 1280
rect 253090 800 253202 1280
rect 254272 0 254384 1280
rect 255454 0 255566 1280
rect 256636 800 256748 1280
rect 257818 0 257930 1280
rect 259000 0 259112 1280
rect 260182 800 260294 1280
rect 261364 0 261476 1280
rect 262546 0 262658 1280
rect 263728 800 263840 1280
rect 264910 0 265022 1280
rect 266092 0 266204 1280
rect 267274 800 267386 1280
rect 268456 0 268568 1280
rect 269638 1175 269752 1280
rect 269638 0 269750 1175
rect 270820 800 270932 1280
rect 272002 0 272114 1280
rect 273184 0 273296 1280
rect 274366 800 274478 1280
rect 275548 0 275660 1280
rect 276730 0 276842 1280
rect 277912 800 278024 1280
rect 279094 0 279206 1280
rect 280276 0 280388 1280
rect 281458 800 281570 1280
rect 282640 0 282752 1280
rect 283822 0 283934 1280
rect 285004 800 285116 1280
rect 286186 0 286298 1280
rect 287368 0 287480 1280
rect 288550 800 288662 1280
rect 289732 0 289844 1280
rect 290914 0 291026 1280
rect 292096 800 292208 1280
rect 293278 0 293390 1280
rect 294460 0 294572 1280
rect 295642 800 295754 1280
rect 296824 0 296936 1280
rect 298006 0 298118 1280
rect 299188 800 299300 1280
rect 300370 0 300482 1280
rect 301552 0 301664 1280
rect 302734 800 302846 1280
rect 303916 0 304028 1280
rect 305098 0 305210 1280
rect 306280 800 306392 1280
rect 307462 0 307574 1280
rect 308644 0 308756 1280
rect 309826 800 309938 1280
rect 311008 0 311120 1280
rect 312190 0 312302 1280
rect 313372 800 313484 1280
rect 314554 0 314666 1280
rect 315736 0 315848 1280
rect 316918 800 317030 1280
rect 318100 0 318212 1280
rect 319282 0 319394 1280
rect 320464 800 320576 1280
rect 321646 0 321758 1280
rect 322828 0 322940 1280
rect 324010 800 324122 1280
rect 325192 0 325304 1280
rect 326374 0 326486 1280
rect 327556 800 327668 1280
rect 328738 0 328850 1280
rect 331102 800 331214 1280
rect 332284 0 332396 1280
rect 333466 0 333578 1280
rect 334648 800 334760 1280
rect 335830 0 335942 1280
rect 338194 800 338306 1280
rect 339376 0 339488 1280
rect 340558 0 340670 1280
rect 341740 800 341852 1280
rect 342922 0 343034 1280
rect 345286 800 345398 1280
rect 346468 0 346580 1280
rect 347650 0 347762 1280
rect 348832 800 348944 1280
rect 350014 0 350126 1280
rect 351196 0 351308 1280
rect 352378 800 352490 1280
rect 353560 0 353672 1280
rect 354742 0 354854 1280
rect 355924 800 356036 1280
rect 357106 0 357218 1280
rect 358288 0 358400 1280
rect 359470 800 359582 1280
rect 360652 0 360764 1280
rect 363016 800 363128 1280
rect 364198 0 364310 1280
rect 365380 0 365492 1280
rect 366562 800 366674 1280
rect 367744 0 367856 1280
rect 370108 800 370220 1280
rect 371290 0 371402 1280
rect 372472 0 372584 1280
rect 373654 800 373766 1280
rect 374836 0 374948 1280
rect 377200 800 377312 1280
rect 378382 0 378494 1280
rect 379564 0 379676 1280
rect 380746 800 380858 1280
rect 381928 0 382040 1280
rect 384292 800 384404 1280
rect 385474 0 385586 1280
rect 386656 0 386768 1280
rect 387838 800 387950 1280
rect 389020 0 389132 1280
rect 391384 800 391496 1280
rect 392566 0 392678 1280
rect 393748 0 393860 1280
rect 394930 800 395042 1280
rect 396112 0 396224 1280
rect 398476 800 398588 1280
rect 399658 0 399770 1280
rect 400840 0 400952 1280
rect 402022 800 402134 1280
rect 403204 0 403316 1280
rect 404386 0 404498 1280
rect 405568 800 405680 1280
rect 406750 0 406862 1280
rect 407932 0 408044 1280
rect 409114 800 409226 1280
rect 410296 0 410408 1280
rect 411478 0 411590 1280
rect 412660 800 412772 1280
rect 413842 0 413954 1280
rect 415024 0 415136 1280
rect 416206 800 416318 1280
rect 417388 0 417500 1280
rect 418570 0 418682 1280
rect 419752 800 419864 1280
rect 420934 0 421046 1280
rect 422116 0 422228 1280
rect 423298 800 423410 1280
rect 424480 0 424592 1280
rect 425662 0 425774 1280
rect 426844 800 426956 1280
rect 428023 1176 428138 1296
rect 431556 1280 431676 6353
rect 458295 5617 458412 412283
rect 435107 5500 458412 5617
rect 458587 412900 458704 412934
rect 435107 1280 435224 5500
rect 458587 4993 458704 412283
rect 438657 4876 458704 4993
rect 458893 412900 459010 412937
rect 438657 1280 438774 4876
rect 458893 4549 459010 412283
rect 442206 4432 459010 4549
rect 459229 412900 459346 412930
rect 442206 1296 442323 4432
rect 459229 3958 459346 412283
rect 445756 3841 459346 3958
rect 459597 412900 459714 412930
rect 445756 1296 445873 3841
rect 459597 3448 459714 412283
rect 460146 412912 460350 412936
rect 547144 412928 547393 413369
rect 552551 412928 559324 413369
rect 460146 412264 460174 412912
rect 460328 412264 460350 412912
rect 466206 412763 473703 412769
rect 466196 412620 559318 412763
rect 466196 412320 466355 412620
rect 460146 412236 460350 412264
rect 460196 16196 460290 412236
rect 466206 410038 466355 412320
rect 473541 412320 559318 412620
rect 473541 410038 473703 412320
rect 466206 409865 473703 410038
rect 580930 369269 581274 369297
rect 580930 367739 580964 369269
rect 581233 367739 581274 369269
rect 580930 367703 581274 367739
rect 582908 368196 583306 368262
rect 580981 367266 581227 367703
rect 580981 366233 581227 366286
rect 582908 365988 582944 368196
rect 583273 365988 583306 368196
rect 582908 365319 583306 365988
rect 580109 361187 581287 361243
rect 580109 360563 580208 361187
rect 581211 360563 581287 361187
rect 583575 361027 584320 361051
rect 583575 360769 583603 361027
rect 584293 360769 584320 361027
rect 583575 360746 584320 360769
rect 580109 360507 581287 360563
rect 577423 356547 577733 357068
rect 577413 356505 577736 356547
rect 577413 355566 577440 356505
rect 577713 355566 577736 356505
rect 577413 355534 577736 355566
rect 577874 353396 577994 357159
rect 578171 356545 578457 357047
rect 578158 356507 578481 356545
rect 578158 355568 578188 356507
rect 578461 355568 578481 356507
rect 578158 355532 578481 355568
rect 580975 355293 581243 355312
rect 580975 354384 581001 355293
rect 581227 354384 581243 355293
rect 580975 354358 581243 354384
rect 577874 353276 580899 353396
rect 567090 316809 568186 316873
rect 567090 315844 567177 316809
rect 568123 316556 568186 316809
rect 568123 316328 573167 316556
rect 568123 315844 568186 316328
rect 567090 315777 568186 315844
rect 569251 315568 570067 315681
rect 569251 314111 569330 315568
rect 569965 314111 570067 315568
rect 569251 313992 570067 314111
rect 571015 314309 572629 314379
rect 571015 313895 571103 314309
rect 572537 313895 572629 314309
rect 571015 313812 572629 313895
rect 571839 311837 573546 311870
rect 571839 311649 571913 311837
rect 573518 311649 573546 311837
rect 571839 311590 573546 311649
rect 571886 311272 573200 311356
rect 512756 283816 513108 283828
rect 512756 283710 512768 283816
rect 513094 283797 513108 283816
rect 513094 283733 515870 283797
rect 513094 283710 513108 283733
rect 512756 283698 513108 283710
rect 511200 279727 511828 279740
rect 511200 279615 511217 279727
rect 511805 279712 511828 279727
rect 511805 279648 516228 279712
rect 511805 279615 511828 279648
rect 511200 279597 511828 279615
rect 513183 268320 513645 268345
rect 513183 268319 515887 268320
rect 513183 268240 513211 268319
rect 513617 268254 515887 268319
rect 513617 268240 513645 268254
rect 513183 268214 513645 268240
rect 515135 267901 515496 267915
rect 515135 267817 515155 267901
rect 515474 267893 515496 267901
rect 515474 267827 516259 267893
rect 515474 267817 515496 267827
rect 515135 267799 515496 267817
rect 514748 267252 515114 267265
rect 514748 267164 514769 267252
rect 515094 267236 515114 267252
rect 515094 267172 516253 267236
rect 515094 267164 515114 267172
rect 514748 267150 515114 267164
rect 513592 265842 514054 265864
rect 513592 265763 513617 265842
rect 514023 265814 514054 265842
rect 514023 265763 515955 265814
rect 513592 265754 515955 265763
rect 513592 265733 514054 265754
rect 514119 265326 514439 265329
rect 514113 265269 514129 265326
rect 514430 265269 516226 265326
rect 514113 265266 516226 265269
rect 460715 264687 515868 264747
rect 460160 16174 460330 16196
rect 460160 15816 460182 16174
rect 460314 15816 460330 16174
rect 460160 15792 460330 15816
rect 449306 3331 459714 3448
rect 449306 1296 449423 3331
rect 460715 3020 460805 264687
rect 452867 2930 460805 3020
rect 461215 264187 515903 264247
rect 428026 0 428138 1176
rect 429208 0 429320 1176
rect 430390 800 430502 1280
rect 431556 1111 431684 1280
rect 431572 0 431684 1111
rect 432754 0 432866 1280
rect 433936 800 434048 1280
rect 435107 1014 435230 1280
rect 435118 0 435230 1014
rect 436300 0 436412 1280
rect 437482 800 437594 1280
rect 438657 981 438776 1280
rect 438664 0 438776 981
rect 439846 0 439958 1280
rect 441028 800 441140 1280
rect 442206 1014 442322 1296
rect 442210 0 442322 1014
rect 443392 0 443504 1014
rect 444574 800 444686 1280
rect 445756 0 445868 1296
rect 449306 1280 449414 1296
rect 452867 1280 452957 2930
rect 461215 2626 461305 264187
rect 510625 263833 510994 263863
rect 510625 263789 510659 263833
rect 456399 2536 461305 2626
rect 461673 263729 510659 263789
rect 456399 1280 456489 2536
rect 461673 2156 461763 263729
rect 510625 263690 510659 263729
rect 510959 263690 510994 263833
rect 510625 263663 510994 263690
rect 511805 263831 512174 263855
rect 511805 263688 511832 263831
rect 512132 263789 512174 263831
rect 512132 263729 516231 263789
rect 512132 263688 512174 263729
rect 511805 263655 512174 263688
rect 513221 260060 513312 260074
rect 513221 259670 513234 260060
rect 513296 259670 513312 260060
rect 513221 259654 513312 259670
rect 513617 260060 513708 260074
rect 513617 259670 513633 260060
rect 513695 259670 513708 260060
rect 513617 259654 513708 259670
rect 514235 259869 514312 259881
rect 463137 248118 463221 249486
rect 463537 248416 463621 249486
rect 463937 248738 464021 249486
rect 464337 249039 464421 249486
rect 464737 249302 464821 249486
rect 464631 249290 464905 249302
rect 464631 249183 464650 249290
rect 464889 249183 464905 249290
rect 464631 249171 464905 249183
rect 464214 249029 464488 249039
rect 464214 248922 464233 249029
rect 464472 248922 464488 249029
rect 464214 248908 464488 248922
rect 463827 248729 464101 248738
rect 463827 248622 463847 248729
rect 464086 248622 464101 248729
rect 463827 248607 464101 248622
rect 463410 248403 463684 248416
rect 463410 248296 463426 248403
rect 463665 248296 463684 248403
rect 463410 248285 463684 248296
rect 463033 248106 463307 248118
rect 463033 247999 463049 248106
rect 463288 247999 463307 248106
rect 463033 247987 463307 247999
rect 463137 2259 463221 247987
rect 463537 2594 463621 248285
rect 463937 2902 464021 248607
rect 464337 3237 464421 248908
rect 464737 3583 464821 249171
rect 513232 238811 513301 259654
rect 513631 239059 513700 259654
rect 514235 259571 514236 259869
rect 514235 246302 514312 259571
rect 529244 249837 529360 249859
rect 523676 249802 523762 249819
rect 523676 249471 523682 249802
rect 523754 249471 523762 249802
rect 523676 249455 523762 249471
rect 523678 246663 523755 249455
rect 529244 249315 529267 249837
rect 529341 249315 529360 249837
rect 529244 249285 529360 249315
rect 529274 247456 529337 249285
rect 571886 248484 571970 311272
rect 573143 310129 573456 311150
rect 573143 310108 573457 310129
rect 573143 309638 573174 310108
rect 573428 309638 573457 310108
rect 573143 309614 573457 309638
rect 580779 273260 580899 353276
rect 582578 314662 583714 314710
rect 582578 314328 582644 314662
rect 583666 314328 583714 314662
rect 582578 314280 583714 314328
rect 562840 248400 571970 248484
rect 577874 273140 580899 273260
rect 529248 247427 529364 247456
rect 529248 246905 529270 247427
rect 529344 246905 529364 247427
rect 529248 246882 529364 246905
rect 523678 246586 562326 246663
rect 514235 246225 561965 246302
rect 561566 245568 561706 245592
rect 561566 244946 561592 245568
rect 561676 244946 561706 245568
rect 561566 244917 561706 244946
rect 513493 239049 513891 239059
rect 513493 238965 513513 239049
rect 513867 238965 513891 239049
rect 513493 238945 513891 238965
rect 513631 238943 513700 238945
rect 513059 238798 513448 238811
rect 513059 238722 513087 238798
rect 513424 238722 513448 238798
rect 513059 238703 513448 238722
rect 513232 238701 513301 238703
rect 516952 168076 517370 168088
rect 516952 167978 516964 168076
rect 517356 168051 517370 168076
rect 517356 167999 521368 168051
rect 517356 167978 517370 167999
rect 516952 167966 517370 167978
rect 517032 163836 517475 163845
rect 517032 163746 517043 163836
rect 517464 163828 517475 163836
rect 517464 163764 521352 163828
rect 517464 163746 517475 163764
rect 517032 163736 517475 163746
rect 475632 133510 538106 133520
rect 475632 133452 537879 133510
rect 538076 133452 538106 133510
rect 475632 133445 538106 133452
rect 475632 3867 475707 133445
rect 475832 133312 538106 133320
rect 475832 133254 536151 133312
rect 536348 133254 538106 133312
rect 475832 133245 538106 133254
rect 475832 4126 475907 133245
rect 476032 133110 538106 133120
rect 476032 133052 534348 133110
rect 534545 133052 538106 133110
rect 476032 133045 538106 133052
rect 476032 4395 476107 133045
rect 476232 132912 538106 132920
rect 476232 132854 534096 132912
rect 534293 132854 538106 132912
rect 476232 132845 538106 132854
rect 476232 4692 476307 132845
rect 476432 132711 538106 132720
rect 476432 132653 533808 132711
rect 534005 132653 538106 132711
rect 476432 132645 538106 132653
rect 476432 4922 476507 132645
rect 476632 132510 538106 132520
rect 476632 132452 533528 132510
rect 533725 132452 538106 132510
rect 476632 132445 538106 132452
rect 476632 5182 476707 132445
rect 511588 78174 512103 78188
rect 511588 77972 511606 78174
rect 512088 78143 512103 78174
rect 512088 78079 516226 78143
rect 512088 77972 512103 78079
rect 511588 77954 512103 77972
rect 511540 74171 512094 74186
rect 511540 74031 511558 74171
rect 512077 74143 512094 74171
rect 512077 74079 516444 74143
rect 512077 74031 512094 74079
rect 511540 74016 512094 74031
rect 513539 62082 516237 62134
rect 513539 46321 513591 62082
rect 513842 61732 516250 61788
rect 513842 47227 513898 61732
rect 514200 56714 516137 56742
rect 513831 47212 513909 47227
rect 513831 46976 513838 47212
rect 513899 46976 513909 47212
rect 513831 46966 513909 46976
rect 513521 46308 513621 46321
rect 513521 46055 513539 46308
rect 513603 46055 513621 46308
rect 513521 46036 513621 46055
rect 514200 45774 514228 56714
rect 514795 56070 516130 56098
rect 478882 45746 514228 45774
rect 478882 5422 478940 45746
rect 514796 45565 514824 56070
rect 479091 45537 514824 45565
rect 515096 50274 516142 50302
rect 479091 5652 479149 45537
rect 515096 45377 515124 50274
rect 515337 47220 515415 47235
rect 515337 46984 515344 47220
rect 515405 46984 515415 47220
rect 515337 46974 515415 46984
rect 479279 45349 515124 45377
rect 479279 5892 479337 45349
rect 515351 45345 515390 46974
rect 560829 45357 561153 45372
rect 560829 45345 560845 45357
rect 515351 45306 560845 45345
rect 560829 45301 560845 45306
rect 561136 45301 561153 45357
rect 560829 45289 561153 45301
rect 479525 45124 534315 45131
rect 479525 45065 534097 45124
rect 534304 45065 534315 45124
rect 479525 45055 534315 45065
rect 479525 6217 479601 45055
rect 479725 44922 534315 44931
rect 479725 44863 533511 44922
rect 533718 44863 534315 44922
rect 479725 44855 534315 44863
rect 479725 6417 479801 44855
rect 479925 44723 534315 44731
rect 479925 44664 531429 44723
rect 531636 44664 534315 44723
rect 479925 44655 534315 44664
rect 479925 6617 480001 44655
rect 480125 44523 534315 44531
rect 480125 44464 531124 44523
rect 531331 44464 534315 44523
rect 480125 44455 534315 44464
rect 480125 6817 480201 44455
rect 480325 44323 534315 44331
rect 480325 44264 530771 44323
rect 530978 44264 534315 44323
rect 480325 44255 534315 44264
rect 480325 7017 480401 44255
rect 480525 44123 534315 44131
rect 480525 44064 526989 44123
rect 527196 44064 534315 44123
rect 480525 44055 534315 44064
rect 480525 7217 480601 44055
rect 480725 43923 534315 43931
rect 480725 43864 525627 43923
rect 525834 43864 534315 43923
rect 480725 43855 534315 43864
rect 480725 7417 480801 43855
rect 480925 43723 534315 43731
rect 480925 43664 523599 43723
rect 523806 43664 534315 43723
rect 480925 43655 534315 43664
rect 480925 7617 481001 43655
rect 522988 43452 523334 43472
rect 522988 43386 522999 43452
rect 523317 43446 523334 43452
rect 523317 43386 561400 43446
rect 522988 43370 561400 43386
rect 561323 9110 561400 43370
rect 542704 9033 561400 9110
rect 480925 7541 538044 7617
rect 480725 7341 534503 7417
rect 480525 7141 530943 7217
rect 480325 6941 527402 7017
rect 480125 6741 523870 6817
rect 479925 6541 520319 6617
rect 479725 6341 516768 6417
rect 479525 6141 513218 6217
rect 479279 5834 509677 5892
rect 479091 5594 506126 5652
rect 478882 5364 502566 5422
rect 476632 5107 499033 5182
rect 476432 4847 495482 4922
rect 476232 4617 491941 4692
rect 476032 4320 488371 4395
rect 475832 4051 484849 4126
rect 475632 3792 481308 3867
rect 464737 3499 477771 3583
rect 464337 3153 474221 3237
rect 463937 2818 470670 2902
rect 463537 2510 467129 2594
rect 463137 2175 463578 2259
rect 459950 2066 461763 2156
rect 459950 1280 460040 2066
rect 463494 1280 463578 2175
rect 467045 1280 467129 2510
rect 470586 1280 470670 2818
rect 474137 1280 474221 3153
rect 477687 1280 477771 3499
rect 481233 1280 481308 3792
rect 484774 1280 484849 4051
rect 488296 1280 488371 4320
rect 491866 1280 491941 4617
rect 495407 1280 495482 4847
rect 498958 1280 499033 5107
rect 502508 1280 502566 5364
rect 506068 1280 506126 5594
rect 509619 1280 509677 5834
rect 513142 1280 513218 6141
rect 516692 1280 516768 6341
rect 520243 1280 520319 6541
rect 523794 1280 523870 6741
rect 527326 1280 527402 6941
rect 530867 1280 530943 7141
rect 534427 1280 534503 7341
rect 537968 1280 538044 7541
rect 542704 1280 542781 9033
rect 561612 8859 561689 244917
rect 545073 8782 561689 8859
rect 545073 1280 545150 8782
rect 561888 8446 561965 246225
rect 549786 8369 561965 8446
rect 549786 1280 549863 8369
rect 562249 8102 562326 246586
rect 553344 8025 562326 8102
rect 553344 1280 553421 8025
rect 562840 7569 562924 248400
rect 577874 247844 577994 273140
rect 578786 272103 579326 272134
rect 578786 272101 579726 272103
rect 578786 271811 578848 272101
rect 579290 271871 579726 272101
rect 579290 271811 579326 271871
rect 578786 271784 579326 271811
rect 578267 270783 579168 270845
rect 578267 270535 578316 270783
rect 579119 270535 579168 270783
rect 578267 270495 579168 270535
rect 583850 270272 584276 270316
rect 583850 269860 583912 270272
rect 584220 269860 584276 270272
rect 578265 269758 579153 269826
rect 583850 269812 584276 269860
rect 578265 269456 578330 269758
rect 579103 269456 579153 269758
rect 578265 269412 579153 269456
rect 579005 267379 579830 267422
rect 579005 267185 579061 267379
rect 579777 267185 579830 267379
rect 579005 267142 579830 267185
rect 555704 7485 562924 7569
rect 563238 247724 577994 247844
rect 578604 266814 579583 266888
rect 555704 1280 555788 7485
rect 563238 7086 563358 247724
rect 563638 246063 563778 246087
rect 563638 245441 563664 246063
rect 563748 245971 563778 246063
rect 578604 245971 578678 266814
rect 579511 266070 579857 266682
rect 579506 266043 579859 266070
rect 579506 265637 579525 266043
rect 579842 265637 579859 266043
rect 579506 265610 579859 265637
rect 563748 245897 578678 245971
rect 563748 245441 563778 245897
rect 563638 245412 563778 245441
rect 566612 239361 566668 239365
rect 566559 239344 566963 239361
rect 566559 239273 566586 239344
rect 566941 239273 566963 239344
rect 566559 239258 566963 239273
rect 566315 239056 566371 239061
rect 566132 239038 566536 239056
rect 566132 238967 566159 239038
rect 566514 238967 566536 239038
rect 566132 238953 566536 238967
rect 565947 238804 566003 238807
rect 565775 238785 566179 238804
rect 565775 238714 565800 238785
rect 566155 238714 566179 238785
rect 565775 238701 566179 238714
rect 565947 80246 566003 238701
rect 566315 80614 566371 238953
rect 566612 80911 566668 239258
rect 566612 80855 580509 80911
rect 566315 80558 580212 80614
rect 565947 80190 579844 80246
rect 579433 42523 579551 42545
rect 579433 42199 579450 42523
rect 579522 42199 579551 42523
rect 579433 42173 579551 42199
rect 579104 42026 579222 42048
rect 579104 41702 579123 42026
rect 579195 41702 579222 42026
rect 579104 41676 579222 41702
rect 579143 26894 579199 41676
rect 579449 26897 579505 42173
rect 579788 26898 579844 80190
rect 579118 26872 579240 26894
rect 579118 26514 579140 26872
rect 579213 26514 579240 26872
rect 579118 26494 579240 26514
rect 579421 26871 579543 26897
rect 579421 26513 579438 26871
rect 579511 26513 579543 26871
rect 579421 26497 579543 26513
rect 579750 26872 579872 26898
rect 580156 26897 580212 80558
rect 580453 26900 580509 80855
rect 582047 27953 583234 27996
rect 582047 27654 582111 27953
rect 583186 27654 583234 27953
rect 582047 27606 583234 27654
rect 579750 26514 579770 26872
rect 579843 26514 579872 26872
rect 579750 26498 579872 26514
rect 580115 26872 580237 26897
rect 580115 26514 580133 26872
rect 580206 26514 580237 26872
rect 580115 26497 580237 26514
rect 580420 26879 580542 26900
rect 580420 26521 580440 26879
rect 580513 26521 580542 26879
rect 580420 26500 580542 26521
rect 582968 25125 583171 27606
rect 582968 24613 583000 25125
rect 583140 24613 583171 25125
rect 582968 20364 583171 24613
rect 582968 19852 582991 20364
rect 583131 19852 583171 20364
rect 563626 15898 563756 15912
rect 563626 15502 563640 15898
rect 563748 15502 563756 15898
rect 563626 15478 563756 15502
rect 582968 15647 583171 19852
rect 559223 6966 563358 7086
rect 446938 0 447050 1063
rect 448120 800 448232 1280
rect 449302 0 449414 1280
rect 450484 0 450596 1096
rect 451666 800 451778 1280
rect 452848 0 452960 1280
rect 454030 0 454142 1280
rect 455212 800 455324 1280
rect 456394 0 456506 1280
rect 457576 1190 457696 1280
rect 457576 0 457688 1190
rect 458758 800 458870 1280
rect 459940 0 460052 1280
rect 461122 0 461234 1280
rect 462304 800 462416 1280
rect 463486 0 463598 1280
rect 464668 1094 464787 1280
rect 464668 0 464780 1094
rect 465850 800 465962 1280
rect 467032 0 467144 1280
rect 468214 1163 468329 1280
rect 468214 0 468326 1163
rect 469396 800 469508 1280
rect 470578 0 470690 1280
rect 471760 0 471872 1280
rect 472942 800 473054 1280
rect 474124 0 474236 1280
rect 475306 0 475418 1280
rect 476488 800 476600 1280
rect 477670 0 477782 1280
rect 478852 0 478964 1280
rect 480034 800 480146 1280
rect 481216 0 481328 1280
rect 482398 0 482510 1280
rect 483580 800 483692 1280
rect 484762 0 484874 1280
rect 485944 0 486056 1280
rect 487126 800 487238 1280
rect 488296 1124 488420 1280
rect 488308 0 488420 1124
rect 489490 0 489602 1280
rect 490672 800 490784 1280
rect 491854 0 491966 1280
rect 493036 0 493148 1280
rect 494218 800 494330 1280
rect 495400 0 495512 1280
rect 496582 0 496694 1280
rect 497764 800 497876 1280
rect 498946 0 499058 1280
rect 500128 0 500240 1280
rect 501310 800 501422 1280
rect 502492 0 502604 1280
rect 503674 0 503786 1280
rect 504856 800 504968 1280
rect 506038 0 506150 1280
rect 507220 0 507332 1280
rect 508402 800 508514 1280
rect 509584 0 509696 1280
rect 510766 0 510878 1280
rect 511948 800 512060 1280
rect 513130 0 513242 1280
rect 514312 0 514424 1280
rect 515494 800 515606 1280
rect 516676 0 516788 1280
rect 517858 0 517970 1280
rect 519040 800 519152 1280
rect 520222 0 520334 1280
rect 521404 0 521516 1280
rect 522586 800 522698 1280
rect 523768 0 523880 1280
rect 524950 0 525062 1280
rect 526132 800 526244 1280
rect 527314 0 527426 1280
rect 528496 0 528608 1280
rect 529678 800 529790 1280
rect 530860 0 530972 1280
rect 532042 0 532154 1280
rect 533224 800 533336 1280
rect 534406 0 534518 1280
rect 535588 0 535700 1280
rect 536770 800 536882 1280
rect 537952 0 538064 1280
rect 539134 0 539246 1280
rect 540316 800 540428 1280
rect 540340 0 540428 800
rect 541498 0 541610 1280
rect 542680 0 542792 1280
rect 543862 800 543974 1280
rect 545044 0 545156 1280
rect 546226 0 546338 1280
rect 547408 800 547520 1280
rect 547422 0 547520 800
rect 548590 0 548702 1280
rect 549772 0 549884 1280
rect 550954 800 551066 1280
rect 550980 0 551066 800
rect 552136 0 552248 1280
rect 553318 0 553430 1280
rect 554500 800 554612 1280
rect 555682 0 555794 1280
rect 556864 0 556976 1280
rect 558046 800 558158 1280
rect 559223 1124 559343 6966
rect 563640 3148 563716 15478
rect 563906 15198 564046 15216
rect 563906 14808 563932 15198
rect 564020 14808 564046 15198
rect 563906 14778 564046 14808
rect 582968 15135 583004 15647
rect 583144 15135 583171 15647
rect 563932 3616 564010 14778
rect 582968 10963 583171 15135
rect 582968 10933 583181 10963
rect 569644 10676 569964 10692
rect 569644 10590 569672 10676
rect 569944 10590 569964 10676
rect 569644 10574 569964 10590
rect 563932 3525 566423 3616
rect 562798 3072 563716 3148
rect 559228 0 559340 1124
rect 560410 0 560522 1445
rect 562798 1280 562874 3072
rect 566345 1280 566423 3525
rect 569868 1280 569946 10574
rect 582968 10421 583002 10933
rect 583142 10421 583181 10933
rect 582968 10391 583181 10421
rect 582968 6190 583171 10391
rect 582968 5664 583003 6190
rect 583137 5664 583171 6190
rect 582968 3856 583171 5664
rect 561592 800 561704 1280
rect 562774 0 562886 1280
rect 563956 0 564068 1280
rect 565138 800 565250 1280
rect 566320 0 566432 1280
rect 567502 0 567614 1280
rect 568684 800 568796 1280
rect 569866 0 569978 1280
rect 571048 0 571160 1280
rect 572230 800 572342 1280
rect 573412 0 573524 1280
rect 574594 0 574706 1280
rect 575776 800 575888 1280
rect 576958 0 577070 1280
rect 578140 0 578252 1280
rect 579322 800 579434 1280
rect 580504 800 580616 1280
rect 581686 800 581798 1280
rect 582868 800 582980 1280
rect 584050 800 584162 1280
<< via2 >>
rect 263662 653984 265591 654713
rect 321200 653975 323129 654704
rect 245788 652377 247717 653106
rect 339074 652368 341003 653097
rect 263662 563984 265591 564713
rect 245788 562377 247717 563106
rect 28395 486659 38334 492430
rect 6256 470365 12269 475393
rect 2262 468578 2494 469256
rect 7494 469100 8300 469236
rect 15660 469083 15889 469755
rect 18241 478121 18645 479537
rect 136929 480414 140755 481050
rect 128886 479271 132750 479922
rect 7523 461352 8290 461984
rect 5436 455115 6072 456528
rect 136913 457377 140759 458053
rect 128913 456233 132752 456791
rect 129000 446760 132676 448269
rect 6459 436151 6743 436988
rect 13424 434895 14366 436724
rect 136929 433457 140750 434133
rect 128909 432251 132750 432842
rect 6378 429877 7086 430832
rect 11697 427828 13585 428240
rect 4522 425868 4717 426541
rect 8126 384475 9182 384757
rect 8553 382858 9115 383290
rect 1730 382608 2548 382780
rect 8241 381897 9368 382289
rect 7617 379740 9223 379992
rect 7609 378984 9228 379239
rect 59802 358268 60356 359034
rect 4993 344467 5879 344582
rect 1564 339376 2527 339574
rect 4983 339220 5982 339653
rect 6789 334800 7923 335356
rect 4974 334263 5809 334449
rect 3091 311780 3736 314581
rect 8496 335696 9359 336159
rect 5395 301251 6315 301415
rect 1959 296191 2922 296389
rect 5290 296044 6335 296534
rect 7102 291597 8352 292119
rect 5396 291105 6049 291271
rect 8908 292471 9750 293051
rect 8301 287438 8561 288005
rect 9412 286596 9675 287240
rect 9050 285653 9285 286322
rect 11839 302797 12083 302878
rect 11835 302596 12079 302677
rect 10745 88436 11391 89075
rect 12471 88436 13117 89075
rect 9045 84367 9901 85362
rect 3580 44203 4529 44764
rect 1484 38894 1684 39496
rect 5712 38923 6434 39422
rect 9153 35396 9363 35996
rect 60381 34422 60444 34705
rect 9132 33660 9845 33908
rect 8266 33163 8753 33376
rect 9136 32419 9849 32667
rect 7258 27214 7592 28409
rect 60541 34422 60604 34705
rect 60701 34422 60764 34705
rect 60861 34422 60924 34705
rect 61021 34422 61084 34705
rect 61181 34422 61244 34705
rect 61341 34422 61404 34705
rect 61501 34422 61564 34705
rect 65259 34421 65322 34661
rect 65419 34421 65482 34661
rect 65579 34421 65642 34661
rect 65739 34421 65802 34661
rect 65899 34421 65962 34661
rect 66059 34421 66122 34661
rect 66219 34421 66282 34661
rect 66379 34421 66442 34661
rect 263662 476584 265591 477313
rect 245788 472377 247717 473106
rect 263662 383984 265591 384713
rect 245788 382377 247717 383106
rect 263662 293984 265591 294713
rect 245788 292377 247717 293106
rect 263662 203984 265591 204713
rect 245788 202377 247717 203106
rect 263662 113984 265591 114713
rect 245788 112377 247717 113106
rect 181967 14869 182409 14965
rect 181554 7340 182266 7436
rect 280236 11032 280439 11088
rect 279888 10904 280091 10960
rect 279573 10776 279722 10832
rect 279262 10648 279398 10704
rect 278859 10521 279049 10577
rect 278570 10391 278691 10447
rect 278154 10263 278357 10319
rect 275217 10135 275420 10191
rect 271663 10009 271866 10065
rect 268139 9881 268342 9937
rect 264562 9751 264765 9807
rect 261017 9624 261220 9680
rect 286531 281121 286590 281299
rect 298623 281046 298693 281284
rect 286731 280434 286790 280629
rect 286931 279306 286990 279501
rect 287131 277218 287190 277413
rect 287331 275123 287390 275318
rect 287531 273032 287590 273227
rect 287731 269860 287790 270055
rect 287931 264595 287990 264802
rect 298423 264095 298493 264296
rect 298223 207988 298293 208190
rect 288131 197431 288190 197629
rect 298023 155388 298093 155592
rect 297823 102891 297893 103096
rect 288309 87051 288390 87253
rect 290122 30361 290933 30905
rect 288835 11032 289038 11088
rect 288461 10904 288664 10960
rect 288257 10776 288460 10832
rect 288062 10648 288265 10704
rect 287865 10520 288068 10576
rect 287663 10392 287866 10448
rect 287464 10264 287667 10320
rect 287255 10137 287458 10193
rect 287069 10008 287272 10064
rect 286866 9880 287069 9936
rect 286679 9752 286882 9808
rect 286461 9624 286664 9680
rect 297359 10474 297562 10530
rect 297555 10346 297758 10402
rect 297753 10218 297956 10274
rect 297960 10089 298163 10145
rect 298158 9962 298361 10018
rect 298354 9834 298557 9890
rect 298894 56610 298962 57142
rect 298896 10620 299168 10678
rect 298550 9706 298753 9762
rect 444372 614087 448011 617699
rect 513911 593259 520276 609778
rect 568944 588943 569285 589315
rect 583568 588859 583746 589372
rect 573573 585613 574366 586727
rect 583874 584260 584212 584564
rect 577145 583409 577661 584173
rect 510907 570179 518330 576926
rect 321200 563975 323129 564704
rect 339074 562368 341003 563097
rect 452351 563112 455990 566724
rect 560571 564711 562698 565066
rect 438947 561526 439446 561647
rect 565447 581487 565813 581852
rect 439355 560950 439854 561071
rect 568964 580566 569295 580907
rect 422782 558790 423705 558959
rect 576075 496743 576616 498421
rect 575013 495447 575808 496291
rect 576790 493993 577757 494849
rect 583490 494882 584168 495102
rect 578317 492070 579412 492276
rect 460200 491736 460638 491840
rect 578266 491321 579420 491568
rect 321200 473975 323129 474704
rect 339074 472368 341003 473097
rect 557782 434769 557961 435818
rect 583321 433815 583433 434170
rect 583313 431416 583425 431771
rect 419509 422017 421145 422228
rect 452329 420650 456074 421269
rect 444386 418708 447969 419339
rect 321200 383975 323129 384704
rect 339074 382368 341003 383097
rect 339074 294368 341003 295097
rect 321212 292187 323141 292916
rect 439388 216140 439512 216572
rect 321200 203975 323129 204704
rect 339074 202368 341003 203097
rect 321200 113975 323129 114704
rect 339074 112368 341003 113097
rect 456314 14942 456522 15732
rect 403156 10474 403359 10530
rect 406710 10346 406913 10402
rect 410268 10218 410471 10274
rect 413816 10088 414019 10144
rect 417353 9961 417556 10017
rect 420889 9832 421092 9888
rect 424463 9705 424666 9761
rect 554002 415181 554622 415365
rect 556144 415189 556764 415373
rect 554002 414441 554622 414625
rect 556144 414449 556764 414633
rect 458295 412283 458412 412900
rect 458587 412283 458704 412900
rect 458893 412283 459010 412900
rect 459229 412283 459346 412900
rect 459597 412283 459714 412900
rect 547393 412928 552551 413369
rect 460174 412264 460328 412912
rect 466355 410038 473541 412620
rect 580964 367739 581233 369269
rect 582944 365988 583273 368196
rect 580208 360563 581211 361187
rect 583603 360769 584293 361027
rect 577440 355566 577713 356505
rect 578188 355568 578461 356507
rect 581001 354384 581227 355293
rect 567177 315844 568123 316809
rect 569330 314111 569965 315568
rect 571103 313895 572537 314309
rect 571913 311649 573518 311837
rect 512768 283710 513094 283816
rect 511217 279615 511805 279727
rect 513211 268240 513617 268319
rect 515155 267817 515474 267901
rect 514769 267164 515094 267252
rect 513617 265763 514023 265842
rect 514129 265269 514430 265326
rect 460182 15816 460314 16174
rect 510659 263690 510959 263833
rect 511832 263688 512132 263831
rect 513234 259670 513296 260060
rect 513633 259670 513695 260060
rect 464650 249183 464889 249290
rect 464233 248922 464472 249029
rect 463847 248622 464086 248729
rect 463426 248296 463665 248403
rect 463049 247999 463288 248106
rect 514236 259571 514312 259869
rect 523682 249471 523754 249802
rect 529267 249315 529341 249837
rect 573174 309638 573428 310108
rect 582644 314328 583666 314662
rect 529270 246905 529344 247427
rect 561592 244946 561676 245568
rect 513513 238965 513867 239049
rect 513087 238722 513424 238798
rect 516964 167978 517356 168076
rect 517043 163746 517464 163836
rect 537879 133452 538076 133510
rect 536151 133254 536348 133312
rect 534348 133052 534545 133110
rect 534096 132854 534293 132912
rect 533808 132653 534005 132711
rect 533528 132452 533725 132510
rect 511606 77972 512088 78174
rect 511558 74031 512077 74171
rect 513838 46976 513899 47212
rect 513539 46055 513603 46308
rect 515344 46984 515405 47220
rect 560845 45301 561136 45357
rect 534097 45065 534304 45124
rect 533511 44863 533718 44922
rect 531429 44664 531636 44723
rect 531124 44464 531331 44523
rect 530771 44264 530978 44323
rect 526989 44064 527196 44123
rect 525627 43864 525834 43923
rect 523599 43664 523806 43723
rect 522999 43386 523317 43452
rect 578848 271811 579290 272101
rect 578316 270535 579119 270783
rect 583912 269860 584220 270272
rect 578330 269456 579103 269758
rect 579061 267185 579777 267379
rect 563664 245441 563748 246063
rect 579525 265637 579842 266043
rect 566586 239273 566941 239344
rect 566159 238967 566514 239038
rect 565800 238714 566155 238785
rect 579450 42199 579522 42523
rect 579123 41702 579195 42026
rect 579140 26514 579213 26872
rect 579438 26513 579511 26871
rect 582111 27654 583186 27953
rect 579770 26514 579843 26872
rect 580133 26514 580206 26872
rect 580440 26521 580513 26879
rect 583000 24613 583140 25125
rect 582991 19852 583131 20364
rect 563640 15502 563748 15898
rect 563932 14808 564020 15198
rect 583004 15135 583144 15647
rect 569672 10590 569944 10676
rect 583002 10421 583142 10933
rect 583003 5664 583137 6190
<< metal3 >>
rect 16994 703100 21994 705600
rect 68994 703100 73994 705600
rect 120994 703100 125994 705600
rect 166394 703100 171394 705600
rect 171694 703100 173894 704800
rect 174194 703100 176394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 705600
rect 223394 703100 225594 704800
rect 225894 703100 228094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 325094 703100 327294 704800
rect 327594 703100 329794 704800
rect 330094 703100 335094 705600
rect 414194 703100 419194 705600
rect 466194 703100 471194 705600
rect 18574 687352 19364 703100
rect 71019 691045 71393 703100
rect 71019 690671 117078 691045
rect 18574 686562 105509 687352
rect 0 683312 2500 686042
rect 0 682498 101676 683312
rect 0 681042 2500 682498
rect 0 649314 8531 649442
rect 0 644833 3472 649314
rect 8318 644833 8531 649314
rect 0 644642 8531 644833
rect 800 639260 8531 639442
rect 800 634779 3494 639260
rect 8340 634779 8531 639260
rect 800 634642 8531 634779
rect 0 564868 9296 565042
rect 0 560414 4054 564868
rect 9132 560414 9296 564868
rect 0 560242 9296 560414
rect 800 554880 9296 555042
rect 800 550426 4066 554880
rect 9144 550426 9296 554880
rect 800 550242 9296 550426
rect 0 512330 1280 512442
rect 914 511260 4453 511427
rect 0 511148 13837 511260
rect 914 511054 4453 511148
rect 800 509966 1280 510078
rect 800 508784 1280 508896
rect 0 507602 1280 507714
rect 100862 507674 101676 682498
rect 99670 507328 102794 507674
rect 0 506420 1280 506532
rect 99670 504650 100018 507328
rect 102298 504650 102794 507328
rect 99670 504204 102794 504650
rect 28157 492430 38565 492612
rect 28157 486659 28395 492430
rect 38334 486659 38565 492430
rect 28157 486422 38565 486659
rect 18196 479537 18710 479594
rect 18196 478121 18241 479537
rect 18645 478121 18710 479537
rect 18196 478064 18710 478121
rect 4420 475393 12415 475493
rect 4420 470365 6256 475393
rect 12269 470365 12415 475393
rect 4420 470219 12415 470365
rect 15621 469755 15920 469792
rect 2247 469256 2512 469278
rect 2247 469220 2262 469256
rect 0 469108 838 469220
rect 1168 469108 2262 469220
rect 2247 468578 2262 469108
rect 2494 469013 2512 469256
rect 7459 469236 8334 469270
rect 7459 469100 7494 469236
rect 8300 469220 8334 469236
rect 15621 469220 15660 469755
rect 8300 469108 15660 469220
rect 8300 469100 8334 469108
rect 7459 469073 8334 469100
rect 15621 469083 15660 469108
rect 15889 469083 15920 469755
rect 15621 469053 15920 469083
rect 2494 468578 2511 469013
rect 2247 468557 2511 468578
rect 0 467926 1280 468038
rect 800 466744 1280 466856
rect 800 465562 1280 465674
rect 0 464380 1280 464492
rect 0 463198 1280 463310
rect 7466 461984 8347 462028
rect 7466 461352 7523 461984
rect 8290 461352 8347 461984
rect 7466 461302 8347 461352
rect 5343 456528 6129 456631
rect 5343 455115 5436 456528
rect 6072 455115 6129 456528
rect 5343 455031 6129 455115
rect 43252 452040 45058 452203
rect 43252 443121 43381 452040
rect 44947 443121 45058 452040
rect 104719 448630 105509 686562
rect 103912 448182 106444 448630
rect 103912 446394 104310 448182
rect 106146 446394 106444 448182
rect 103912 446048 106444 446394
rect 6447 436988 6755 437005
rect 6447 436151 6459 436988
rect 6743 436590 6755 436988
rect 13382 436724 14416 436761
rect 6743 436151 12660 436590
rect 6447 436150 12660 436151
rect 6447 436136 6755 436150
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 12220 430688 12660 436150
rect 13382 434895 13424 436724
rect 14366 436708 14416 436724
rect 43252 436708 45058 443121
rect 14366 434902 45058 436708
rect 14366 434895 14416 434902
rect 13382 434848 14416 434895
rect 74070 430688 74510 430689
rect 12220 430248 74510 430688
rect 6302 429814 7162 429877
rect 11637 428240 13660 428297
rect 11637 427828 11697 428240
rect 13585 427828 13660 428240
rect 11637 427782 13660 427828
rect 4484 426541 4759 426575
rect 4484 426125 4522 426541
rect 1061 425998 4522 426125
rect 0 425886 4522 425998
rect 1061 425868 4522 425886
rect 4717 425998 4759 426541
rect 4717 425886 4760 425998
rect 4717 425868 4759 425886
rect 1061 425840 4759 425868
rect 4484 425830 4759 425840
rect 0 424704 1280 424816
rect 800 423522 1280 423634
rect 800 422340 1280 422452
rect 0 421158 1280 421270
rect 0 419976 1280 420088
rect 74070 384820 74510 430248
rect 8087 384757 9234 384793
rect 8087 384475 8126 384757
rect 9182 384475 9234 384757
rect 8087 384441 9234 384475
rect 73769 384777 74673 384820
rect 73769 384033 73831 384777
rect 74622 384033 74673 384777
rect 73769 383978 74673 384033
rect 8490 383290 9178 383354
rect 8490 382858 8553 383290
rect 9115 382858 9178 383290
rect 1694 382780 2576 382812
rect 8490 382807 9178 382858
rect 1694 382776 1730 382780
rect 0 382664 1730 382776
rect 1694 382608 1730 382664
rect 2548 382608 2576 382780
rect 1694 382578 2576 382608
rect 8167 382289 9436 382347
rect 8167 381897 8241 382289
rect 9368 381897 9436 382289
rect 8167 381846 9436 381897
rect 0 381482 1280 381594
rect 800 380300 1280 380412
rect 7571 379992 9262 380019
rect 7571 379740 7617 379992
rect 9223 379740 9262 379992
rect 7571 379709 9262 379740
rect 7566 379239 9272 379263
rect 800 379118 1280 379230
rect 7566 378984 7609 379239
rect 9228 378984 9272 379239
rect 7566 378955 9272 378984
rect 0 377936 2454 378048
rect 1363 376882 2182 376909
rect 1363 376866 1392 376882
rect 0 376754 1288 376866
rect 1353 376754 1392 376866
rect 1363 376729 1392 376754
rect 2159 376729 2182 376882
rect 1363 376706 2182 376729
rect 2342 359856 2454 377936
rect 59760 364712 60412 364756
rect 59760 363848 59828 364712
rect 60326 363848 60412 364712
rect 2342 359756 17556 359856
rect 17456 358678 17556 359756
rect 59760 359034 60412 363848
rect 59760 358268 59802 359034
rect 60356 358268 60412 359034
rect 59760 358208 60412 358268
rect 116704 347944 117078 690671
rect 115878 347766 118262 347944
rect 115878 345626 116072 347766
rect 118072 345626 118262 347766
rect 115878 345460 118262 345626
rect 4957 344582 14018 344626
rect 4957 344467 4993 344582
rect 5879 344467 14018 344582
rect 4957 344428 14018 344467
rect 4935 339653 6035 339688
rect 1528 339574 2590 339613
rect 1528 339554 1564 339574
rect 0 339442 1564 339554
rect 1528 339376 1564 339442
rect 2527 339376 2590 339574
rect 1528 339348 2590 339376
rect 4935 339220 4983 339653
rect 5982 339220 6035 339653
rect 4935 339168 6035 339220
rect 0 338260 1280 338372
rect 800 337078 1280 337190
rect 11107 336581 11768 336620
rect 11107 336225 11146 336581
rect 8442 336159 11146 336225
rect 800 335896 1280 336008
rect 8442 335696 8496 336159
rect 9359 335696 11146 336159
rect 8442 335652 11146 335696
rect 11723 335652 11768 336581
rect 8442 335630 11768 335652
rect 11107 335605 11768 335630
rect 6704 335356 8008 335437
rect 0 334714 1280 334826
rect 6704 334800 6789 335356
rect 7923 334800 8008 335356
rect 6704 334714 8008 334800
rect 4944 334464 7776 334465
rect 4943 334449 7776 334464
rect 4943 334263 4974 334449
rect 5809 334263 7776 334449
rect 4943 334245 7776 334263
rect 4943 334244 5832 334245
rect 0 333532 1280 333644
rect 3032 314581 3801 314651
rect 3032 311780 3091 314581
rect 3736 311780 3801 314581
rect 3032 311699 3801 311780
rect 7556 307000 7776 334245
rect 13820 317188 14018 344428
rect 25656 318928 26056 318962
rect 25656 318190 25702 318928
rect 26022 318190 26056 318928
rect 25656 318140 26056 318190
rect 34316 317188 34516 317838
rect 13820 316988 34516 317188
rect 35156 316348 35356 317838
rect 7556 306618 7588 307000
rect 7747 306618 7776 307000
rect 7556 306587 7776 306618
rect 8577 316148 35356 316348
rect 8577 301432 8775 316148
rect 50006 310650 50498 310690
rect 50006 310072 50036 310650
rect 50460 310072 50498 310650
rect 10005 308203 10187 308217
rect 10005 307782 10019 308203
rect 10174 307782 10187 308203
rect 10005 302786 10187 307782
rect 50006 306986 50498 310072
rect 10005 302398 10018 302786
rect 10174 302398 10187 302786
rect 10005 302386 10187 302398
rect 10647 306338 10847 306354
rect 10647 305956 10668 306338
rect 10827 305956 10847 306338
rect 50006 306142 50036 306986
rect 50462 306142 50498 306986
rect 50006 306104 50498 306142
rect 5372 301415 8775 301432
rect 5372 301251 5395 301415
rect 6315 301251 8775 301415
rect 5372 301234 8775 301251
rect 5194 296534 6467 296612
rect 1917 296389 2979 296430
rect 1917 296332 1959 296389
rect 0 296220 1959 296332
rect 1917 296191 1959 296220
rect 2922 296191 2979 296389
rect 1917 296165 2979 296191
rect 5194 296044 5290 296534
rect 6335 296044 6467 296534
rect 5194 295966 6467 296044
rect 0 295038 1280 295150
rect 800 293856 1280 293968
rect 8863 293051 9807 293093
rect 800 292674 1280 292786
rect 8863 292471 8908 293051
rect 9750 292471 9807 293051
rect 8863 292434 9807 292471
rect 7037 292119 8427 292167
rect 0 291492 1280 291604
rect 7037 291597 7102 292119
rect 8352 291597 8427 292119
rect 7037 291557 8427 291597
rect 5372 291288 6070 291289
rect 10647 291288 10847 305956
rect 11825 302878 12095 302887
rect 11825 302797 11839 302878
rect 12083 302797 12095 302878
rect 11825 302787 12095 302797
rect 11825 302677 12092 302686
rect 11825 302596 11835 302677
rect 12079 302596 12092 302677
rect 11825 302587 12092 302596
rect 5372 291271 10847 291288
rect 5372 291105 5396 291271
rect 6049 291105 10847 291271
rect 5372 291088 10847 291105
rect 0 290310 1280 290422
rect 8280 288005 10428 288028
rect 8280 287438 8301 288005
rect 8561 287991 10428 288005
rect 8561 287438 9820 287991
rect 8280 287428 9820 287438
rect 10389 287428 10428 287991
rect 8280 287404 10428 287428
rect 5195 287240 9698 287259
rect 5195 287221 9412 287240
rect 5195 286612 5242 287221
rect 6400 286612 9412 287221
rect 5195 286596 9412 286612
rect 9675 286596 9698 287240
rect 122792 287156 123728 703100
rect 168369 697685 168783 703100
rect 146740 697271 168783 697685
rect 128832 653097 132832 656117
rect 128832 652362 128918 653097
rect 132733 652362 132832 653097
rect 128832 595370 132832 652362
rect 136832 654723 140832 656662
rect 136832 653988 136910 654723
rect 140725 653988 140832 654723
rect 136832 644370 140832 653988
rect 136832 639691 136986 644370
rect 140674 639691 140832 644370
rect 128823 595069 132844 595370
rect 128823 589599 129074 595069
rect 132598 589599 132844 595069
rect 128823 589258 132844 589599
rect 128832 563093 132832 589258
rect 128832 562358 128910 563093
rect 132725 562358 132832 563093
rect 128832 479922 132832 562358
rect 128832 479271 128886 479922
rect 132750 479271 132832 479922
rect 128832 475246 132832 479271
rect 128832 472150 128924 475246
rect 132768 472150 132832 475246
rect 128832 456791 132832 472150
rect 128832 456233 128913 456791
rect 132752 456233 132832 456791
rect 128832 448269 132832 456233
rect 128832 446760 129000 448269
rect 132676 446760 132832 448269
rect 128832 432842 132832 446760
rect 128832 432251 128909 432842
rect 132750 432251 132832 432842
rect 128832 383136 132832 432251
rect 128832 382381 128923 383136
rect 132755 382381 132832 383136
rect 128832 380144 132832 382381
rect 128832 379827 128918 380144
rect 132762 379827 132832 380144
rect 128832 377026 132832 379827
rect 128832 376582 128962 377026
rect 132722 376582 132832 377026
rect 128832 364692 132832 376582
rect 128832 363838 128893 364692
rect 132628 363838 132832 364692
rect 128832 310649 132832 363838
rect 128832 310102 128934 310649
rect 132738 310102 132832 310649
rect 128832 293105 132832 310102
rect 128832 292378 128935 293105
rect 132733 292378 132832 293105
rect 5195 286568 9698 286596
rect 121856 286830 124852 287156
rect 7775 286322 9309 286351
rect 7775 286306 9050 286322
rect 7775 285650 7809 286306
rect 8396 285653 9050 286306
rect 9285 285653 9309 286322
rect 8396 285650 9309 285653
rect 7775 285616 9309 285650
rect 121856 284192 122182 286830
rect 124562 284192 124852 286830
rect 121856 283880 124852 284192
rect 10297 253568 11453 253569
rect 1102 253310 11453 253568
rect 0 253198 11453 253310
rect 1102 252959 11453 253198
rect 0 252016 1280 252128
rect 800 250834 1280 250946
rect 800 249652 1280 249764
rect 0 248470 1280 248582
rect 0 247288 1280 247400
rect 0 220396 9632 220488
rect 0 215890 4310 220396
rect 9440 215890 9632 220396
rect 10297 220080 11453 252959
rect 10297 220037 11458 220080
rect 10297 218186 10348 220037
rect 10300 218145 10348 218186
rect 11403 218145 11458 220037
rect 10300 218090 11458 218145
rect 0 215688 9632 215890
rect 800 210358 9632 210488
rect 800 205852 4284 210358
rect 9414 205852 9632 210358
rect 800 205688 9632 205852
rect 128832 203118 132832 292378
rect 128832 202363 128929 203118
rect 132761 202363 132832 203118
rect 0 178310 9505 178488
rect 0 173829 3756 178310
rect 8602 173829 9505 178310
rect 0 173688 9505 173829
rect 128832 173511 132832 202363
rect 128832 168834 129023 173511
rect 132621 168834 132832 173511
rect 800 168320 9505 168488
rect 800 163839 3676 168320
rect 8522 163839 9505 168320
rect 800 163688 9505 163839
rect 994 125688 3264 125821
rect 0 125576 3264 125688
rect 994 125450 3264 125576
rect 0 124394 1280 124506
rect 800 123212 1280 123324
rect 800 122030 1280 122142
rect 0 120848 1280 120960
rect 0 119666 1280 119778
rect 2893 98583 3264 125450
rect 118902 117189 124253 117235
rect 118902 116572 122080 117189
rect 124173 116572 124253 117189
rect 118902 116521 124253 116572
rect 118902 115235 119616 116521
rect 15185 114521 119616 115235
rect 8077 113162 10345 113393
rect 15185 113254 15899 114521
rect 8077 109813 8320 113162
rect 10127 110355 10345 113162
rect 128832 113106 132832 168834
rect 128832 112351 128914 113106
rect 132746 112351 132832 113106
rect 10127 109813 10693 110355
rect 8077 109555 10693 109813
rect 4331 107789 6732 108048
rect 4331 104052 4550 107789
rect 6568 104653 6732 107789
rect 6568 104052 10693 104653
rect 4331 103853 10693 104052
rect 4331 103820 6732 103853
rect 2893 98212 10004 98583
rect 2849 95180 9960 95551
rect 2849 82602 3220 95180
rect 984 82466 3220 82602
rect 0 82354 3220 82466
rect 984 82231 3220 82354
rect 5652 92763 9983 93563
rect 5652 83268 6452 92763
rect 7440 91563 9983 92363
rect 7440 85421 8240 91563
rect 7419 85362 11196 85421
rect 7419 85317 9045 85362
rect 9901 85317 11196 85362
rect 7419 84414 7550 85317
rect 11060 84414 11196 85317
rect 7419 84367 9045 84414
rect 9901 84367 11196 84414
rect 7419 84273 11196 84367
rect 5652 83143 9429 83268
rect 5652 82240 5768 83143
rect 9278 82240 9429 83143
rect 5652 82120 9429 82240
rect 0 81172 1280 81284
rect 44761 81065 45051 88677
rect 2863 80775 45051 81065
rect 128832 85335 132832 112351
rect 128832 84353 128916 85335
rect 132725 84353 132832 85335
rect 800 79990 1280 80102
rect 800 78808 1280 78920
rect 0 77626 1280 77738
rect 0 76444 1280 76556
rect 2863 45952 3153 80775
rect 3859 79506 4961 79573
rect 3859 78534 3917 79506
rect 4887 78781 4961 79506
rect 4887 78538 4962 78781
rect 4887 78534 4961 78538
rect 2063 45722 3154 45952
rect 2063 45662 3153 45722
rect 1456 39496 1714 39528
rect 1456 39244 1484 39496
rect 0 39132 1484 39244
rect 1456 38894 1484 39132
rect 1684 38894 1714 39496
rect 1456 38866 1714 38894
rect 0 37950 1280 38062
rect 800 36768 1280 36880
rect 800 35586 1280 35698
rect 2063 34609 2353 45662
rect 3859 44867 4961 78534
rect 3503 44764 4961 44867
rect 3503 44203 3580 44764
rect 4529 44226 4961 44764
rect 128832 56959 132832 84353
rect 128832 53284 128967 56959
rect 132708 53284 132832 56959
rect 4529 44203 4633 44226
rect 3503 44125 4633 44203
rect 5652 39422 6511 39493
rect 5652 38923 5712 39422
rect 6434 38923 6511 39422
rect 5652 38883 6511 38923
rect 9094 35996 9417 36046
rect 9094 35396 9153 35996
rect 9363 35396 9417 35996
rect 9094 35350 9417 35396
rect 1092 34516 2353 34609
rect 0 34404 2353 34516
rect 1092 34319 2353 34404
rect 9103 33954 9409 35350
rect 60376 34705 60456 42355
rect 60376 34422 60381 34705
rect 60444 34422 60456 34705
rect 60376 34413 60456 34422
rect 60536 34705 60616 42355
rect 60536 34422 60541 34705
rect 60604 34422 60616 34705
rect 60536 34413 60616 34422
rect 60696 34705 60776 42355
rect 60696 34422 60701 34705
rect 60764 34422 60776 34705
rect 60696 34413 60776 34422
rect 60856 34705 60936 42355
rect 60856 34422 60861 34705
rect 60924 34422 60936 34705
rect 60856 34413 60936 34422
rect 61016 34705 61096 42355
rect 61016 34422 61021 34705
rect 61084 34422 61096 34705
rect 61016 34413 61096 34422
rect 61176 34705 61256 42355
rect 61176 34422 61181 34705
rect 61244 34422 61256 34705
rect 61176 34413 61256 34422
rect 61336 34705 61416 42355
rect 61336 34422 61341 34705
rect 61404 34422 61416 34705
rect 61336 34413 61416 34422
rect 61496 34705 61576 42355
rect 61496 34422 61501 34705
rect 61564 34422 61576 34705
rect 61496 34413 61576 34422
rect 65252 34661 65332 42355
rect 65252 34421 65259 34661
rect 65322 34421 65332 34661
rect 65252 34413 65332 34421
rect 65412 34661 65492 42355
rect 65412 34421 65419 34661
rect 65482 34421 65492 34661
rect 65412 34413 65492 34421
rect 65572 34661 65652 42355
rect 65572 34421 65579 34661
rect 65642 34421 65652 34661
rect 65572 34413 65652 34421
rect 65732 34661 65812 42355
rect 65732 34421 65739 34661
rect 65802 34421 65812 34661
rect 65732 34413 65812 34421
rect 65892 34661 65972 42355
rect 65892 34421 65899 34661
rect 65962 34421 65972 34661
rect 65892 34413 65972 34421
rect 66052 34661 66132 42355
rect 66052 34421 66059 34661
rect 66122 34421 66132 34661
rect 66052 34413 66132 34421
rect 66212 34661 66292 42355
rect 66212 34421 66219 34661
rect 66282 34421 66292 34661
rect 66212 34413 66292 34421
rect 66372 34661 66452 42355
rect 66372 34421 66379 34661
rect 66442 34421 66452 34661
rect 66372 34413 66452 34421
rect 9065 33908 9908 33954
rect 9065 33660 9132 33908
rect 9845 33660 9908 33908
rect 9065 33610 9908 33660
rect 128832 33416 132832 53284
rect 1131 33334 1444 33416
rect 0 33222 1444 33334
rect 1131 33126 1444 33222
rect 1626 33376 132832 33416
rect 1626 33163 8266 33376
rect 8753 33163 132832 33376
rect 1626 33126 132832 33163
rect 9061 32667 119190 32718
rect 9061 32419 9136 32667
rect 9849 32468 119190 32667
rect 9849 32419 113278 32468
rect 9061 32376 113278 32419
rect 9069 32373 9912 32376
rect 113034 31500 113278 32376
rect 118898 31500 119190 32468
rect 113034 31270 119190 31500
rect 128832 28804 132832 33126
rect 136832 564708 140832 639691
rect 136832 563973 136911 564708
rect 140726 563973 140832 564708
rect 136832 481050 140832 563973
rect 136832 480414 136929 481050
rect 140755 480414 140832 481050
rect 136832 477303 140832 480414
rect 136832 476568 136918 477303
rect 140733 476568 140832 477303
rect 136832 458053 140832 476568
rect 136832 457377 136913 458053
rect 140759 457377 140832 458053
rect 136832 434133 140832 457377
rect 136832 433457 136929 434133
rect 140750 433457 140832 434133
rect 136832 401010 140832 433457
rect 136832 391475 137099 401010
rect 140611 391475 140832 401010
rect 136832 384711 140832 391475
rect 136832 383956 136941 384711
rect 140773 383956 140832 384711
rect 136832 379269 140832 383956
rect 136832 378850 136999 379269
rect 140729 378850 140832 379269
rect 136832 362468 140832 378850
rect 136832 361328 136912 362468
rect 140668 361328 140832 362468
rect 136832 309624 140832 361328
rect 136832 309106 136918 309624
rect 140746 309106 140832 309624
rect 136832 294706 140832 309106
rect 136832 293979 136946 294706
rect 140744 293979 140832 294706
rect 136832 204723 140832 293979
rect 136832 203968 136923 204723
rect 140755 203968 140832 204723
rect 136832 114737 140832 203968
rect 146740 146616 147154 697271
rect 220111 693525 220373 703100
rect 160762 693263 220373 693525
rect 145758 146268 148578 146616
rect 145758 143960 146008 146268
rect 148318 143960 148578 146268
rect 145758 143656 148578 143960
rect 136832 113982 136938 114737
rect 140770 113982 140832 114737
rect 136832 83186 140832 113982
rect 136832 82204 136942 83186
rect 140751 82204 140832 83186
rect 136832 40865 140832 82204
rect 160762 66334 161024 693263
rect 331404 680832 331796 703100
rect 415856 686754 416308 703100
rect 467586 686834 468038 703100
rect 511394 698944 516194 705600
rect 511394 693868 511510 698944
rect 516020 693868 516194 698944
rect 511394 693672 516194 693868
rect 521394 698932 526194 705600
rect 567394 703100 572394 705600
rect 521394 693856 521554 698932
rect 526064 693856 526194 698932
rect 521394 693672 526194 693856
rect 415856 686302 427878 686754
rect 331404 680440 424246 680832
rect 263426 654713 265741 654863
rect 263426 653984 263662 654713
rect 265591 653984 265741 654713
rect 263426 653791 265741 653984
rect 321050 654704 323365 654854
rect 321050 653975 321200 654704
rect 323129 653975 323365 654704
rect 321050 653782 323365 653975
rect 245574 653106 247889 653256
rect 245574 652377 245788 653106
rect 247717 652377 247889 653106
rect 245574 652184 247889 652377
rect 338902 653097 341217 653247
rect 338902 652368 339074 653097
rect 341003 652368 341217 653097
rect 338902 652175 341217 652368
rect 423854 607278 424246 680440
rect 422464 606998 426030 607278
rect 422464 604042 422844 606998
rect 425668 604042 426030 606998
rect 422464 603712 426030 604042
rect 283206 567908 284412 567940
rect 283206 567566 283246 567908
rect 284368 567566 284412 567908
rect 283206 567534 284412 567566
rect 263426 564713 265741 564863
rect 263426 563984 263662 564713
rect 265591 563984 265741 564713
rect 263426 563791 265741 563984
rect 245574 563106 247889 563256
rect 245574 562377 245788 563106
rect 247717 562377 247889 563106
rect 245574 562184 247889 562377
rect 263426 477313 265741 477463
rect 263426 476584 263662 477313
rect 265591 476584 265741 477313
rect 263426 476391 265741 476584
rect 245574 473106 247889 473256
rect 245574 472377 245788 473106
rect 247717 472377 247889 473106
rect 245574 472184 247889 472377
rect 263426 384713 265741 384863
rect 263426 383984 263662 384713
rect 265591 383984 265741 384713
rect 263426 383791 265741 383984
rect 245574 383106 247889 383256
rect 245574 382377 245788 383106
rect 247717 382377 247889 383106
rect 245574 382184 247889 382377
rect 283377 296533 283739 567534
rect 321050 564704 323365 564854
rect 321050 563975 321200 564704
rect 323129 563975 323365 564704
rect 321050 563782 323365 563975
rect 338902 563097 341217 563247
rect 338902 562368 339074 563097
rect 341003 562368 341217 563097
rect 338902 562175 341217 562368
rect 422747 558994 422879 558998
rect 422745 558959 423751 558994
rect 422745 558790 422782 558959
rect 423705 558790 423751 558959
rect 422745 558762 423751 558790
rect 284377 478603 284838 478643
rect 284377 477428 284414 478603
rect 284791 477428 284838 478603
rect 284377 477375 284838 477428
rect 282617 296171 283739 296533
rect 263426 294713 265741 294863
rect 263426 293984 263662 294713
rect 265591 293984 265741 294713
rect 263426 293791 265741 293984
rect 245574 293106 247889 293256
rect 245574 292377 245788 293106
rect 247717 292377 247889 293106
rect 245574 292184 247889 292377
rect 282617 265845 282979 296171
rect 283533 295162 283999 295188
rect 283533 293605 283572 295162
rect 283964 293605 283999 295162
rect 283533 293564 283999 293605
rect 283579 271101 283937 293564
rect 284417 280007 284775 477375
rect 321050 474704 323365 474854
rect 321050 473975 321200 474704
rect 323129 473975 323365 474704
rect 321050 473782 323365 473975
rect 338902 473097 341217 473247
rect 338902 472368 339074 473097
rect 341003 472368 341217 473097
rect 338902 472175 341217 472368
rect 419480 422228 421176 422253
rect 419480 422017 419509 422228
rect 421145 422017 421176 422228
rect 419480 421993 421176 422017
rect 419623 387551 419844 421993
rect 285445 387330 419844 387551
rect 285445 280317 285684 387330
rect 285962 386083 287206 386139
rect 285962 385971 286018 386083
rect 285957 385768 286018 385971
rect 287145 385768 287206 386083
rect 285957 385713 287206 385768
rect 285957 281005 286200 385713
rect 321050 384704 323365 384854
rect 321050 383975 321200 384704
rect 323129 383975 323365 384704
rect 321050 383782 323365 383975
rect 338902 383097 341217 383247
rect 338902 382368 339074 383097
rect 341003 382368 341217 383097
rect 338902 382175 341217 382368
rect 338902 295097 341217 295247
rect 338902 294368 339074 295097
rect 341003 294368 341217 295097
rect 338902 294175 341217 294368
rect 321062 292916 323377 293065
rect 321062 292187 321212 292916
rect 323141 292187 323377 292916
rect 422747 292556 422879 558762
rect 423789 499585 424196 499588
rect 423770 499533 424448 499585
rect 423770 497872 423834 499533
rect 424381 497872 424448 499533
rect 423770 497813 424448 497872
rect 423789 293301 424196 497813
rect 427426 430644 427878 686302
rect 430574 686382 468038 686834
rect 426340 430286 428862 430644
rect 426340 428204 426592 430286
rect 428498 428204 428862 430286
rect 426340 427878 428862 428204
rect 321062 291994 323377 292187
rect 421275 292454 422940 292556
rect 421275 292005 421370 292454
rect 422855 292005 422940 292454
rect 421275 291915 422940 292005
rect 423790 291985 424196 293301
rect 423790 291865 425460 291985
rect 423790 291416 423897 291865
rect 425382 291416 425460 291865
rect 423790 291344 425460 291416
rect 423790 291343 423933 291344
rect 289080 288800 290237 288826
rect 289080 288789 302955 288800
rect 289080 288524 289130 288789
rect 290210 288552 302955 288789
rect 290210 288524 290237 288552
rect 289080 288488 290237 288524
rect 289072 287319 290229 287341
rect 289072 287302 302388 287319
rect 289072 287037 289114 287302
rect 290194 287071 302388 287302
rect 290194 287037 290229 287071
rect 289072 287003 290229 287037
rect 289065 286661 290222 286695
rect 289065 286396 289110 286661
rect 290190 286643 290222 286661
rect 290190 286396 301839 286643
rect 289065 286395 301839 286396
rect 289065 286357 290222 286395
rect 299307 285969 299931 286011
rect 299307 285048 299365 285969
rect 299882 285813 299931 285969
rect 300260 285959 300884 286012
rect 300260 285834 300312 285959
rect 299882 285048 299932 285813
rect 299307 284990 299932 285048
rect 286495 281299 288828 281308
rect 286495 281121 286531 281299
rect 286590 281121 288828 281299
rect 297766 281284 298736 281292
rect 297766 281158 298623 281284
rect 286495 281109 288828 281121
rect 298586 281046 298623 281158
rect 298693 281046 298736 281284
rect 298586 281038 298736 281046
rect 285957 280762 288872 281005
rect 297697 280768 298234 280973
rect 298029 280721 298234 280768
rect 299727 280721 299932 284990
rect 286670 280629 288877 280641
rect 286670 280434 286731 280629
rect 286790 280434 288877 280629
rect 298029 280516 299932 280721
rect 300259 285038 300312 285834
rect 300829 285038 300884 285959
rect 300259 284991 300884 285038
rect 286670 280420 288877 280434
rect 285445 280078 288869 280317
rect 284417 279649 288988 280007
rect 286876 279501 288851 279515
rect 286876 279306 286931 279501
rect 286990 279306 288851 279501
rect 286876 279294 288851 279306
rect 284759 278775 285073 278813
rect 284759 278144 284796 278775
rect 285034 278455 285073 278775
rect 285034 278144 288988 278455
rect 284759 278097 288988 278144
rect 284759 278096 285073 278097
rect 287075 277413 288857 277423
rect 287075 277218 287131 277413
rect 287190 277218 288857 277413
rect 287075 277202 288857 277218
rect 285142 276685 285477 276725
rect 285142 276044 285179 276685
rect 285438 276363 285477 276685
rect 285438 276044 288988 276363
rect 285142 276005 288988 276044
rect 285142 276002 285477 276005
rect 287288 275318 288937 275331
rect 287288 275123 287331 275318
rect 287390 275123 288937 275318
rect 287288 275110 288937 275123
rect 285646 274532 285965 274561
rect 285646 273948 285676 274532
rect 285943 274271 285965 274532
rect 285943 273948 288988 274271
rect 285646 273913 288988 273948
rect 285646 273912 285965 273913
rect 287474 273227 288851 273239
rect 287474 273032 287531 273227
rect 287590 273032 288851 273227
rect 287474 273018 288851 273032
rect 283579 270743 288988 271101
rect 287713 270055 288851 270069
rect 287713 269860 287731 270055
rect 287790 269860 288851 270055
rect 287713 269848 288851 269860
rect 282617 265483 288992 265845
rect 300259 265342 300621 284991
rect 297732 264980 300621 265342
rect 287918 264802 288850 264809
rect 287918 264595 287931 264802
rect 287990 264595 288850 264802
rect 287918 264588 288850 264595
rect 297873 264296 298534 264306
rect 297873 264095 298423 264296
rect 298493 264095 298534 264296
rect 297873 264085 298534 264095
rect 297732 208872 299585 209234
rect 297873 208190 298325 208198
rect 297873 207988 298223 208190
rect 298293 207988 298325 208190
rect 297873 207977 298325 207988
rect 301591 207217 301839 286395
rect 302140 207766 302388 287071
rect 302707 208333 302955 288552
rect 427838 287992 428290 287995
rect 430574 287992 431026 686382
rect 467586 686276 468038 686382
rect 568648 683460 569100 703100
rect 433826 683008 569100 683460
rect 426826 287604 431158 287992
rect 426826 284006 427136 287604
rect 430734 284006 431158 287604
rect 426826 283660 431158 284006
rect 433826 211589 434278 683008
rect 583100 680372 585600 683784
rect 436838 679920 585600 680372
rect 433802 211499 434337 211589
rect 436838 211581 437290 679920
rect 583100 678784 585600 679920
rect 444177 654693 448177 655482
rect 444177 653958 444265 654693
rect 448080 653958 448177 654693
rect 444177 640383 448177 653958
rect 444177 635697 444374 640383
rect 448011 635697 448177 640383
rect 444177 617699 448177 635697
rect 444177 614087 444372 617699
rect 448011 614087 448177 617699
rect 444177 564713 448177 614087
rect 444177 563978 444283 564713
rect 448098 563978 448177 564713
rect 438929 561647 439466 561660
rect 438929 561526 438947 561647
rect 439446 561526 439466 561647
rect 438929 561509 439466 561526
rect 438977 386935 439077 561509
rect 439337 561071 439874 561084
rect 439337 560950 439355 561071
rect 439854 560950 439874 561071
rect 439337 560933 439874 560950
rect 438962 386918 439091 386935
rect 438962 386616 438977 386918
rect 439074 386616 439091 386918
rect 438962 386597 439091 386616
rect 439385 216600 439485 560933
rect 444177 491676 448177 563978
rect 452177 653093 456177 655103
rect 452177 652358 452277 653093
rect 456092 652358 456177 653093
rect 452177 566724 456177 652358
rect 573658 645170 584800 645384
rect 573658 640732 573828 645170
rect 578952 640732 584800 645170
rect 573658 640584 584800 640732
rect 573658 635200 585600 635384
rect 573658 630762 573842 635200
rect 578966 630762 585600 635200
rect 573658 630584 585600 630762
rect 513415 609778 520733 610315
rect 508780 595050 510602 595116
rect 513415 595070 513911 609778
rect 508780 594750 508882 595050
rect 510528 594964 510602 595050
rect 510528 594750 510602 594800
rect 508780 594670 510602 594750
rect 513414 594741 513911 595070
rect 509568 592207 509766 594670
rect 513415 593259 513911 594741
rect 520276 593259 520733 609778
rect 513415 592789 520733 593259
rect 520989 594964 521187 594969
rect 520989 594800 546963 594964
rect 520989 592207 521187 594800
rect 546799 593848 546963 594800
rect 509568 592009 521187 592207
rect 565682 590272 583582 590384
rect 583722 590272 585600 590384
rect 565682 581897 565794 590272
rect 583556 589372 583758 589415
rect 568861 589315 569347 589367
rect 568861 588943 568944 589315
rect 569285 588943 569347 589315
rect 568861 588870 569347 588943
rect 565411 581852 565859 581897
rect 565411 581487 565447 581852
rect 565813 581487 565859 581852
rect 510422 576926 518844 577547
rect 510422 570179 510907 576926
rect 518330 570179 518844 576926
rect 510422 569612 518844 570179
rect 452177 563112 452351 566724
rect 455990 563112 456177 566724
rect 452177 563094 456177 563112
rect 452177 562359 452281 563094
rect 456096 562359 456177 563094
rect 452177 500973 456177 562359
rect 549766 558443 549932 573064
rect 452177 500838 452220 500973
rect 456132 500838 456177 500973
rect 452177 492443 456177 500838
rect 458275 558277 549932 558443
rect 452154 492374 456203 492443
rect 452154 491981 452284 492374
rect 456101 491981 456203 492374
rect 452154 491916 456203 491981
rect 444177 491240 444298 491676
rect 448085 491240 448177 491676
rect 444177 474702 448177 491240
rect 444177 473967 444287 474702
rect 448102 473967 448177 474702
rect 444177 419339 448177 473967
rect 444177 418708 444386 419339
rect 447969 418708 448177 419339
rect 444177 384710 448177 418708
rect 444177 383975 444261 384710
rect 448076 383975 448177 384710
rect 444177 356155 448177 383975
rect 444177 355510 444363 356155
rect 448074 355510 448177 356155
rect 440097 355012 440420 355040
rect 440097 354020 440123 355012
rect 440396 354020 440420 355012
rect 440097 292569 440420 354020
rect 444177 310336 448177 355510
rect 444177 309389 444353 310336
rect 448020 309389 448177 310336
rect 444177 298680 448177 309389
rect 444174 298616 448177 298680
rect 444174 297698 444258 298616
rect 448110 297698 448177 298616
rect 444174 297624 448177 297698
rect 444177 296686 448177 297624
rect 444177 295951 444240 296686
rect 448055 295951 448177 296686
rect 440097 292246 443003 292569
rect 442680 277338 443003 292246
rect 442680 277307 443004 277338
rect 442680 276714 442709 277307
rect 442977 276714 443004 277307
rect 442680 276686 443004 276714
rect 440905 274403 441261 274429
rect 440905 273577 440930 274403
rect 441236 273577 441261 274403
rect 440905 273540 441261 273577
rect 439358 216572 439534 216600
rect 439358 216140 439388 216572
rect 439512 216140 439534 216572
rect 439358 216120 439534 216140
rect 433802 209657 433885 211499
rect 434271 209657 434337 211499
rect 433802 209517 434337 209657
rect 436812 211474 437347 211581
rect 436812 209632 436894 211474
rect 437280 209632 437347 211474
rect 436812 209509 437347 209632
rect 440954 208333 441202 273540
rect 302707 208085 441202 208333
rect 302140 207518 441168 207766
rect 301591 206969 440418 207217
rect 433807 206427 434337 206497
rect 164205 206339 165944 206388
rect 164205 205964 164278 206339
rect 165881 206326 165944 206339
rect 165881 205964 284977 206326
rect 164205 205915 165944 205964
rect 263426 204713 265741 204863
rect 263426 203984 263662 204713
rect 265591 203984 265741 204713
rect 263426 203791 265741 203984
rect 245574 203106 247889 203256
rect 245574 202377 245788 203106
rect 247717 202377 247889 203106
rect 245574 202184 247889 202377
rect 284615 198677 284977 205964
rect 423098 205978 425103 206052
rect 423098 205913 423193 205978
rect 335855 205551 423193 205913
rect 321050 204704 323365 204854
rect 321050 203975 321200 204704
rect 323129 203975 323365 204704
rect 321050 203782 323365 203975
rect 335855 203068 336217 205551
rect 423098 205481 423193 205551
rect 424985 205481 425103 205978
rect 423098 205407 425103 205481
rect 433807 204374 433860 206427
rect 434276 205863 434337 206427
rect 436810 206411 437341 206501
rect 434276 204374 434338 205863
rect 433807 204288 434338 204374
rect 436810 204358 436868 206411
rect 437284 204358 437341 206411
rect 436810 204292 437341 204358
rect 338902 203097 341217 203247
rect 335855 202913 336216 203068
rect 302702 202551 336216 202913
rect 284615 198315 288992 198677
rect 288080 197629 288851 197641
rect 288080 197431 288131 197629
rect 288190 197431 288851 197629
rect 288080 197420 288851 197431
rect 302702 156634 303064 202551
rect 338902 202368 339074 203097
rect 341003 202368 341217 203097
rect 338902 202175 341217 202368
rect 423369 196209 424989 196278
rect 423369 195753 423476 196209
rect 424871 195753 424989 196209
rect 423369 195667 424989 195753
rect 297732 156272 303064 156634
rect 297691 155592 298110 155598
rect 297691 155388 298023 155592
rect 298093 155388 298110 155592
rect 297691 155377 298110 155388
rect 164488 117154 166291 117229
rect 164488 116604 164579 117154
rect 166211 117050 166291 117154
rect 423929 117077 424144 195667
rect 433855 167330 434271 204288
rect 431050 167041 434772 167330
rect 431050 163637 431353 167041
rect 434495 163637 434772 167041
rect 431050 163361 434772 163637
rect 166211 116688 284809 117050
rect 166211 116604 166291 116688
rect 164488 116525 166291 116604
rect 263426 114713 265741 114863
rect 263426 113984 263662 114713
rect 265591 113984 265741 114713
rect 263426 113791 265741 113984
rect 245574 113106 247889 113256
rect 245574 112377 245788 113106
rect 247717 112377 247889 113106
rect 245574 112184 247889 112377
rect 284447 88283 284809 116688
rect 301275 116862 424144 117077
rect 297734 103780 299642 104142
rect 284447 87921 288992 88283
rect 288275 87253 288851 87263
rect 288275 87051 288309 87253
rect 288390 87051 288851 87253
rect 288275 87042 288851 87051
rect 159752 66158 162288 66334
rect 159752 63802 159964 66158
rect 162104 63802 162288 66158
rect 159752 63598 162288 63802
rect 298862 57142 298998 57176
rect 298862 56798 298894 57142
rect 297852 56610 298894 56798
rect 298962 56798 298998 57142
rect 298962 56610 299006 56798
rect 297852 56577 299006 56610
rect 301275 47122 301490 116862
rect 321050 114704 323365 114854
rect 321050 113975 321200 114704
rect 323129 113975 323365 114704
rect 321050 113782 323365 113975
rect 338902 113097 341217 113247
rect 338902 112368 339074 113097
rect 341003 112368 341217 113097
rect 338902 112175 341217 112368
rect 436856 68598 437272 204292
rect 440170 74427 440418 206969
rect 440920 156125 441168 207518
rect 440920 155284 440954 156125
rect 441137 155284 441168 156125
rect 440920 155233 441168 155284
rect 442680 156796 443003 276686
rect 442680 156171 442705 156796
rect 442983 156171 443003 156796
rect 442680 78961 443003 156171
rect 444177 202455 448177 295951
rect 444177 201720 444285 202455
rect 448100 201720 448177 202455
rect 444177 180774 448177 201720
rect 444177 179958 444303 180774
rect 448071 179958 448177 180774
rect 444177 114711 448177 179958
rect 452177 473120 456177 491916
rect 452177 472385 452283 473120
rect 456098 472385 456177 473120
rect 452177 421269 456177 472385
rect 452177 420650 452329 421269
rect 456074 420650 456177 421269
rect 452177 383127 456177 420650
rect 458275 412900 458441 558277
rect 550058 558151 550224 573064
rect 458275 412283 458295 412900
rect 458412 412283 458441 412900
rect 458275 412236 458441 412283
rect 458567 557985 550224 558151
rect 458567 412900 458733 557985
rect 550363 557846 550529 573064
rect 458567 412283 458587 412900
rect 458704 412283 458733 412900
rect 458567 412236 458733 412283
rect 458872 557680 550529 557846
rect 458872 412900 459038 557680
rect 550698 557511 550864 573064
rect 458872 412283 458893 412900
rect 459010 412283 459038 412900
rect 458872 412236 459038 412283
rect 459207 557345 550864 557511
rect 459207 412900 459373 557345
rect 552764 557145 552972 573064
rect 565411 565115 565859 581487
rect 568985 581000 569244 588870
rect 583556 588859 583568 589372
rect 583746 589202 583758 589372
rect 583746 589090 585600 589202
rect 583746 588859 583758 589090
rect 583556 588790 583758 588859
rect 584320 587908 584800 588020
rect 573463 586727 574467 586813
rect 573463 585613 573573 586727
rect 574366 585613 574467 586727
rect 584320 586726 584800 586838
rect 573463 585534 574467 585613
rect 584320 585544 585600 585656
rect 583830 584564 584262 584602
rect 583830 584260 583874 584564
rect 584212 584474 584262 584564
rect 584212 584362 585600 584474
rect 584212 584260 584262 584362
rect 583830 584232 584262 584260
rect 577087 584173 577726 584230
rect 577087 583409 577145 584173
rect 577661 583409 577726 584173
rect 577087 583360 577726 583409
rect 568892 580907 569368 581000
rect 568892 580566 568964 580907
rect 569295 580566 569368 580907
rect 568892 580524 569368 580566
rect 560525 565066 565859 565115
rect 560525 564711 560571 565066
rect 562698 564711 565859 565066
rect 560525 564667 565859 564711
rect 459207 412283 459229 412900
rect 459346 412283 459373 412900
rect 459207 412236 459373 412283
rect 459573 556937 552972 557145
rect 459573 412900 459781 556937
rect 575498 556038 584800 556162
rect 575498 551600 575644 556038
rect 580768 551600 584800 556038
rect 575498 551362 584800 551600
rect 575498 546004 585600 546162
rect 575498 541566 575630 546004
rect 580754 541566 585600 546004
rect 575498 541362 585600 541566
rect 460880 500977 461847 501013
rect 460880 500842 460928 500977
rect 461800 500962 461847 500977
rect 461800 500850 583574 500962
rect 583714 500850 585600 500962
rect 461800 500842 461847 500850
rect 460880 500810 461847 500842
rect 557755 499780 584508 499829
rect 557755 499668 585600 499780
rect 557755 499598 584508 499668
rect 460166 491840 460662 491858
rect 460166 491736 460200 491840
rect 460638 491736 460662 491840
rect 460166 491710 460662 491736
rect 460176 412936 460318 491710
rect 557755 435818 557986 499598
rect 575990 498421 576687 498523
rect 584320 498486 584800 498598
rect 575990 496743 576075 498421
rect 576616 496743 576687 498421
rect 584320 497304 584800 497416
rect 575990 496650 576687 496743
rect 574914 496291 575907 496393
rect 574914 495447 575013 496291
rect 575808 495447 575907 496291
rect 584320 496122 585600 496234
rect 574914 495358 575907 495447
rect 583438 495102 584234 495148
rect 576700 494849 577862 494922
rect 576700 493993 576790 494849
rect 577757 493993 577862 494849
rect 583438 494882 583490 495102
rect 584168 495052 584234 495102
rect 584168 494940 585600 495052
rect 584168 494882 584234 494940
rect 583438 494838 584234 494882
rect 576700 493929 577862 493993
rect 578266 492276 579461 492320
rect 578266 492070 578317 492276
rect 579412 492070 579461 492276
rect 578266 492032 579461 492070
rect 578225 491568 579451 491594
rect 578225 491321 578266 491568
rect 579420 491321 579451 491568
rect 578225 491282 579451 491321
rect 584320 456428 585600 456540
rect 584320 455246 585600 455358
rect 584320 454064 584800 454176
rect 584320 452882 584800 452994
rect 557755 434769 557782 435818
rect 557961 434769 557986 435818
rect 557755 434744 557986 434769
rect 583321 451700 585600 451812
rect 475894 434151 479604 434328
rect 583321 434178 583433 451700
rect 584320 450518 585600 450630
rect 475894 425383 476138 434151
rect 479384 425383 479604 434151
rect 583313 434170 583443 434178
rect 583313 433815 583321 434170
rect 583433 433815 583443 434170
rect 583313 433801 583443 433815
rect 583321 433794 583433 433801
rect 583313 431779 583425 431796
rect 583305 431771 583434 431779
rect 583305 431416 583313 431771
rect 583425 431416 583434 431771
rect 583305 431407 583434 431416
rect 475894 425155 479604 425383
rect 475901 413650 478420 425155
rect 556073 415400 556847 415414
rect 553923 415373 556852 415400
rect 553923 415365 556144 415373
rect 553923 415181 554002 415365
rect 554622 415189 556144 415365
rect 556764 415189 556852 415373
rect 554622 415181 556852 415189
rect 553923 415150 556852 415181
rect 553923 415145 554697 415150
rect 556073 414660 556847 414674
rect 553923 414633 556852 414660
rect 553923 414625 556144 414633
rect 553923 414441 554002 414625
rect 554622 414449 556144 414625
rect 556764 414449 556852 414633
rect 554622 414441 556852 414449
rect 553923 414410 556852 414441
rect 553923 414405 554697 414410
rect 475901 413369 552664 413650
rect 459573 412283 459597 412900
rect 459714 412283 459781 412900
rect 459573 412236 459781 412283
rect 460146 412912 460350 412936
rect 475901 412928 547393 413369
rect 552551 412928 552664 413369
rect 475901 412913 552664 412928
rect 460146 412264 460174 412912
rect 460328 412264 460350 412912
rect 460146 412236 460350 412264
rect 466206 412620 473703 412769
rect 466206 410038 466355 412620
rect 473541 410038 473703 412620
rect 466206 409865 473703 410038
rect 583313 407390 583425 431407
rect 584320 412006 585600 412118
rect 584320 410824 585600 410936
rect 584320 409642 584800 409754
rect 584320 408460 584800 408572
rect 583313 407278 585600 407390
rect 584320 406096 585600 406208
rect 580563 384575 581315 384602
rect 580563 384268 580603 384575
rect 581287 384268 581315 384575
rect 580563 384240 581315 384268
rect 452177 382392 452289 383127
rect 456104 382392 456177 383127
rect 452177 358012 456177 382392
rect 580951 369297 581251 384240
rect 580930 369269 581274 369297
rect 580930 367739 580964 369269
rect 581233 367739 581274 369269
rect 580930 367703 581274 367739
rect 582908 368196 583306 368262
rect 582908 365988 582944 368196
rect 583273 365988 583306 368196
rect 582908 365946 583306 365988
rect 584320 365584 585600 365696
rect 584320 364402 585600 364514
rect 584320 363220 584800 363332
rect 584320 362038 584800 362150
rect 580109 361187 581287 361243
rect 580109 360563 580208 361187
rect 581211 360563 581287 361187
rect 583575 361027 584320 361051
rect 583575 360769 583603 361027
rect 584293 360968 584320 361027
rect 584293 360856 585600 360968
rect 584293 360769 584320 360856
rect 583575 360746 584320 360769
rect 580109 360507 581287 360563
rect 584320 359674 585600 359786
rect 452177 357386 452253 358012
rect 456061 357386 456177 358012
rect 452177 306969 456177 357386
rect 575087 358018 576450 358087
rect 575087 357360 575167 358018
rect 576400 357954 576450 358018
rect 576400 357952 578452 357954
rect 576400 357413 578492 357952
rect 576400 357360 576450 357413
rect 575087 357299 576450 357360
rect 577413 356505 577736 356547
rect 578162 356545 578492 357413
rect 575056 356137 576386 356209
rect 575056 355501 575129 356137
rect 576287 356099 576386 356137
rect 577413 356099 577440 356505
rect 576287 355566 577440 356099
rect 577713 355566 577736 356505
rect 576287 355539 577736 355566
rect 576287 355501 576386 355539
rect 577413 355534 577736 355539
rect 578158 356534 578492 356545
rect 578158 356507 578481 356534
rect 578158 355568 578188 356507
rect 578461 355568 578481 356507
rect 578158 355532 578481 355568
rect 575056 355432 576386 355501
rect 580975 355293 581243 355312
rect 579047 354648 580446 354683
rect 579047 354641 579107 354648
rect 579038 354393 579107 354641
rect 580386 354641 580446 354648
rect 580975 354641 581001 355293
rect 580386 354393 581001 354641
rect 579038 354384 581001 354393
rect 581227 354384 581243 355293
rect 579038 354373 581243 354384
rect 579047 354363 580446 354373
rect 580975 354358 581243 354373
rect 581417 320362 583522 320474
rect 583662 320362 585600 320474
rect 567090 316809 568186 316873
rect 567090 315844 567177 316809
rect 568123 315844 568186 316809
rect 567090 315777 568186 315844
rect 569251 315568 570067 315681
rect 569251 314111 569330 315568
rect 569965 314111 570067 315568
rect 569251 313992 570067 314111
rect 571015 314309 572629 314379
rect 571015 313895 571103 314309
rect 572537 313895 572629 314309
rect 571015 313812 572629 313895
rect 452177 306064 452287 306969
rect 456063 306064 456177 306969
rect 564294 311870 571876 311874
rect 564294 311837 573546 311870
rect 564294 311649 571913 311837
rect 573518 311649 573546 311837
rect 564294 311590 573546 311649
rect 564294 306535 564578 311590
rect 565520 310201 566349 310311
rect 565520 309073 565640 310201
rect 566219 310131 566349 310201
rect 566219 310129 573438 310131
rect 566219 310108 573457 310129
rect 566219 309638 573174 310108
rect 573428 309638 573457 310108
rect 566219 309614 573457 309638
rect 566219 309612 573438 309614
rect 566219 309073 566349 309612
rect 565520 308923 566349 309073
rect 452177 295119 456177 306064
rect 564207 306470 564666 306535
rect 564207 305360 564258 306470
rect 564610 305360 564666 306470
rect 564207 305306 564666 305360
rect 581417 298437 581529 320362
rect 581836 319292 584444 319299
rect 581836 319180 585600 319292
rect 581836 319179 584444 319180
rect 581398 298423 581537 298437
rect 581398 297880 581414 298423
rect 513455 297785 581414 297880
rect 581521 297785 581537 298423
rect 513455 297768 581537 297785
rect 513455 295800 513567 297768
rect 581398 297765 581537 297768
rect 581836 297452 581956 319179
rect 584320 317998 584800 318110
rect 584320 316816 584800 316928
rect 584320 315746 584383 315747
rect 584320 315634 585600 315746
rect 582578 314662 583714 314710
rect 582578 314328 582644 314662
rect 583666 314564 583714 314662
rect 583666 314452 585600 314564
rect 583666 314328 583714 314452
rect 582578 314280 583714 314328
rect 582324 298422 582463 298444
rect 582324 297784 582339 298422
rect 582446 297784 582463 298422
rect 582324 297772 582463 297784
rect 514759 297332 581956 297452
rect 513239 295774 513783 295800
rect 513239 295445 513273 295774
rect 513751 295445 513783 295774
rect 513239 295414 513783 295445
rect 513455 295410 513567 295414
rect 452177 294384 452291 295119
rect 456106 294384 456177 295119
rect 452177 293534 456177 294384
rect 452177 292590 452238 293534
rect 456120 292590 456177 293534
rect 452177 200344 456177 292590
rect 495026 283932 495434 283962
rect 495026 283618 495054 283932
rect 495406 283828 495434 283932
rect 495406 283816 513108 283828
rect 495406 283710 512768 283816
rect 513094 283710 513108 283816
rect 495406 283698 513108 283710
rect 495406 283618 495434 283698
rect 495026 283590 495434 283618
rect 497587 279858 498079 279892
rect 497587 279505 497633 279858
rect 498017 279741 498079 279858
rect 498017 279727 511828 279741
rect 498017 279615 511217 279727
rect 511805 279615 511828 279727
rect 498017 279597 511828 279615
rect 498017 279505 498079 279597
rect 497587 279457 498079 279505
rect 513183 268319 513645 268345
rect 513183 268240 513211 268319
rect 513617 268240 513645 268319
rect 513183 268214 513645 268240
rect 510621 263833 512179 263855
rect 510621 263690 510659 263833
rect 510959 263831 512179 263833
rect 510959 263690 511832 263831
rect 510621 263688 511832 263690
rect 512132 263688 512179 263831
rect 510621 263663 512179 263688
rect 513231 260074 513304 268214
rect 514759 267265 514879 297332
rect 515159 296932 581956 297052
rect 515159 267915 515279 296932
rect 581836 274880 581956 296932
rect 582337 276052 582449 297772
rect 582337 275940 583756 276052
rect 583896 275940 585600 276052
rect 581836 274870 584437 274880
rect 581836 274760 585600 274870
rect 584320 274758 585600 274760
rect 584320 273576 584800 273688
rect 567084 272396 568176 272468
rect 567084 271604 567218 272396
rect 568058 272131 568176 272396
rect 584320 272394 584800 272506
rect 578786 272131 579326 272134
rect 568058 272101 579327 272131
rect 568058 271811 578848 272101
rect 579290 271811 579327 272101
rect 568058 271784 579327 271811
rect 568058 271604 568176 271784
rect 567084 271516 568176 271604
rect 584320 271212 585600 271324
rect 578267 270783 579168 270845
rect 578267 270535 578316 270783
rect 579119 270535 579168 270783
rect 578267 270495 579168 270535
rect 583850 270272 584276 270316
rect 583850 269860 583912 270272
rect 584220 270142 584276 270272
rect 584220 270030 585600 270142
rect 584220 269860 584276 270030
rect 578265 269758 579153 269826
rect 583850 269812 584276 269860
rect 578265 269456 578330 269758
rect 579103 269456 579153 269758
rect 578265 269412 579153 269456
rect 515135 267901 515496 267915
rect 515135 267817 515155 267901
rect 515474 267817 515496 267901
rect 515135 267799 515496 267817
rect 515159 267798 515279 267799
rect 564129 267662 564765 267696
rect 514748 267252 515114 267265
rect 514748 267164 514769 267252
rect 515094 267164 515114 267252
rect 514748 267150 515114 267164
rect 564129 267178 564172 267662
rect 564723 267417 564765 267662
rect 579005 267417 579830 267422
rect 564723 267379 579830 267417
rect 564723 267185 579061 267379
rect 579777 267185 579830 267379
rect 564723 267178 579830 267185
rect 564129 267142 579830 267178
rect 564129 267137 579030 267142
rect 564129 267136 564765 267137
rect 579506 266066 579859 266070
rect 565523 266043 579859 266066
rect 565523 266037 579525 266043
rect 513592 265842 514054 265864
rect 513592 265763 513617 265842
rect 514023 265763 514054 265842
rect 513592 265733 514054 265763
rect 513626 260074 513699 265733
rect 565523 265643 565565 266037
rect 566309 265643 579525 266037
rect 565523 265637 579525 265643
rect 579842 265637 579859 266043
rect 565523 265617 579859 265637
rect 579506 265610 579859 265617
rect 514120 265329 514440 265335
rect 514119 265326 514440 265329
rect 514119 265269 514129 265326
rect 514430 265269 514440 265326
rect 514119 265266 514440 265269
rect 514120 265258 514440 265266
rect 513221 260060 513312 260074
rect 513221 259670 513234 260060
rect 513296 259670 513312 260060
rect 513221 259654 513312 259670
rect 513617 260060 513708 260074
rect 513617 259670 513633 260060
rect 513695 259670 513708 260060
rect 514237 259883 514310 265258
rect 513617 259654 513708 259670
rect 514227 259869 514319 259883
rect 514227 259571 514236 259869
rect 514312 259571 514319 259869
rect 514227 259554 514319 259571
rect 523696 249819 523756 251445
rect 525056 250820 525116 251453
rect 525004 250793 525194 250820
rect 525004 250571 525018 250793
rect 525156 250571 525194 250793
rect 525004 250533 525194 250571
rect 525056 250518 525116 250533
rect 525001 250059 525191 250090
rect 525001 249837 525018 250059
rect 525156 249837 525191 250059
rect 529267 249859 529327 251494
rect 529595 250610 529655 251443
rect 529531 250576 529721 250610
rect 529991 250601 530051 251435
rect 530330 250614 530390 251435
rect 529531 250354 529560 250576
rect 529698 250354 529721 250576
rect 529531 250323 529721 250354
rect 529915 250560 530105 250601
rect 529915 250338 529935 250560
rect 530073 250338 530105 250560
rect 529915 250314 530105 250338
rect 530275 250584 530465 250614
rect 530275 250362 530303 250584
rect 530441 250362 530465 250584
rect 530275 250327 530465 250362
rect 530330 250324 530390 250327
rect 523676 249802 523762 249819
rect 525001 249803 525191 249837
rect 529244 249837 529360 249859
rect 523676 249471 523682 249802
rect 523754 249471 523762 249802
rect 523676 249455 523762 249471
rect 464631 249290 464905 249302
rect 464631 249256 464650 249290
rect 463016 249196 464650 249256
rect 464631 249183 464650 249196
rect 464889 249256 464905 249290
rect 525056 249256 525116 249803
rect 529244 249315 529267 249837
rect 529341 249315 529360 249837
rect 529529 249788 529719 249827
rect 529529 249566 529549 249788
rect 529687 249566 529719 249788
rect 529529 249540 529719 249566
rect 529911 249795 530101 249833
rect 529911 249573 529940 249795
rect 530078 249573 530101 249795
rect 529911 249546 530101 249573
rect 530275 249808 530465 249849
rect 530275 249586 530288 249808
rect 530426 249586 530465 249808
rect 530275 249562 530465 249586
rect 529244 249285 529360 249315
rect 464889 249196 525116 249256
rect 464889 249183 464905 249196
rect 464631 249171 464905 249183
rect 464214 249029 464488 249039
rect 464214 248994 464233 249029
rect 463010 248934 464233 248994
rect 464214 248922 464233 248934
rect 464472 248994 464488 249029
rect 529595 248994 529655 249540
rect 464472 248934 529655 248994
rect 464472 248922 464488 248934
rect 464214 248908 464488 248922
rect 463827 248729 464101 248738
rect 463827 248710 463847 248729
rect 463020 248650 463847 248710
rect 463827 248622 463847 248650
rect 464086 248710 464101 248729
rect 529991 248710 530051 249546
rect 464086 248650 530051 248710
rect 464086 248622 464101 248650
rect 463827 248607 464101 248622
rect 463410 248403 463684 248416
rect 463410 248385 463426 248403
rect 462999 248325 463426 248385
rect 463410 248296 463426 248325
rect 463665 248385 463684 248403
rect 530330 248385 530390 249562
rect 463665 248325 530390 248385
rect 463665 248296 463684 248325
rect 463410 248285 463684 248296
rect 463033 248106 463307 248118
rect 463033 248092 463049 248106
rect 462945 248028 463049 248092
rect 463033 247999 463049 248028
rect 463288 248092 463307 248106
rect 533205 248092 533269 251445
rect 463288 248028 533269 248092
rect 463288 247999 463307 248028
rect 463033 247987 463307 247999
rect 529248 247427 529364 247456
rect 529248 246905 529270 247427
rect 529344 246905 529364 247427
rect 529248 246882 529364 246905
rect 529285 239336 529345 246882
rect 563638 246063 563778 246087
rect 561566 245568 561706 245592
rect 561566 244946 561592 245568
rect 561676 245552 561706 245568
rect 563638 245552 563664 246063
rect 561676 245467 563664 245552
rect 561676 244946 561706 245467
rect 563638 245441 563664 245467
rect 563748 246047 563778 246063
rect 563748 245962 563779 246047
rect 563748 245441 563778 245962
rect 563638 245412 563778 245441
rect 561566 244917 561706 244946
rect 574794 240690 584800 240830
rect 566559 239344 566963 239361
rect 566559 239336 566586 239344
rect 529285 239276 566586 239336
rect 566559 239273 566586 239276
rect 566941 239273 566963 239344
rect 566559 239258 566963 239273
rect 513493 239051 513891 239059
rect 566132 239051 566536 239056
rect 513493 239049 566538 239051
rect 513493 238965 513513 239049
rect 513867 239038 566538 239049
rect 513867 238967 566159 239038
rect 566514 238967 566538 239038
rect 513867 238965 566538 238967
rect 513493 238962 566538 238965
rect 513493 238945 513891 238962
rect 566132 238953 566536 238962
rect 513059 238802 513448 238811
rect 565775 238802 566179 238804
rect 513059 238798 566184 238802
rect 513059 238722 513087 238798
rect 513424 238785 566184 238798
rect 513424 238722 565800 238785
rect 513059 238714 565800 238722
rect 566155 238714 566184 238785
rect 513059 238713 566184 238714
rect 513059 238703 513448 238713
rect 565775 238701 566179 238713
rect 574794 236252 574934 240690
rect 580058 236252 584800 240690
rect 574794 236030 584800 236252
rect 574794 230660 585600 230830
rect 574794 226222 574962 230660
rect 580086 226222 585600 230660
rect 574794 226030 585600 226222
rect 452177 199609 452266 200344
rect 456081 199609 456177 200344
rect 452177 191899 456177 199609
rect 574794 196850 584800 197030
rect 574794 192412 574896 196850
rect 580020 192412 584800 196850
rect 574794 192230 584800 192412
rect 452177 187251 452333 191899
rect 455990 187251 456177 191899
rect 452177 177590 456177 187251
rect 574794 186806 585600 187030
rect 574794 182368 574908 186806
rect 580032 182368 585600 186806
rect 574794 182230 585600 182368
rect 452176 177478 456177 177590
rect 452176 176624 452276 177478
rect 456058 176624 456177 177478
rect 452176 176524 456177 176624
rect 444177 113976 444260 114711
rect 448075 113976 448177 114711
rect 444177 92247 448177 113976
rect 444177 91356 444290 92247
rect 448055 91356 448177 92247
rect 442643 78912 443060 78961
rect 442643 77894 442690 78912
rect 443023 77894 443060 78912
rect 442643 77852 443060 77894
rect 440169 74403 440421 74427
rect 440169 73811 440192 74403
rect 440394 73811 440421 74403
rect 440169 73781 440421 73811
rect 440170 73739 440418 73781
rect 436838 67677 437290 68598
rect 435826 67289 440158 67677
rect 435826 63691 436136 67289
rect 439734 63691 440158 67289
rect 435826 63345 440158 63691
rect 136832 31547 137083 40865
rect 140503 31547 140832 40865
rect 136832 30160 140832 31547
rect 285697 46840 289043 47069
rect 297617 46907 301490 47122
rect 7204 28409 7656 28442
rect 7204 27214 7258 28409
rect 7592 27214 7656 28409
rect 7204 27149 7656 27214
rect 7353 22229 7582 27149
rect 128832 23480 129020 28804
rect 132614 23480 132832 28804
rect 128832 23252 132832 23480
rect 285697 22229 285926 46840
rect 444177 34284 448177 91356
rect 452177 113100 456177 176524
rect 492899 168076 517370 168088
rect 492899 167978 516964 168076
rect 517356 167978 517370 168076
rect 492899 167966 517370 167978
rect 492899 156356 493021 167966
rect 494548 163836 517475 163845
rect 494548 163746 517043 163836
rect 517464 163746 517475 163836
rect 494548 163736 517475 163746
rect 492646 156342 493210 156356
rect 492646 156162 492662 156342
rect 493194 156162 493210 156342
rect 492646 156148 493210 156162
rect 494548 155756 494657 163736
rect 493979 155736 494657 155756
rect 493979 155582 494004 155736
rect 494639 155582 494657 155736
rect 493979 155562 494657 155582
rect 574794 152256 584800 152430
rect 574794 147818 575156 152256
rect 580280 147818 584800 152256
rect 574794 147630 584800 147818
rect 574794 142194 585600 142430
rect 574794 137756 575102 142194
rect 580226 137756 585600 142194
rect 574794 137630 585600 137756
rect 533287 132161 533347 134543
rect 533603 132520 533663 134443
rect 533885 132720 533945 134443
rect 534169 132920 534229 134443
rect 534417 133120 534477 134443
rect 536217 133320 536281 134443
rect 537953 133520 538017 134443
rect 537870 133510 538083 133520
rect 537870 133452 537879 133510
rect 538076 133452 538083 133510
rect 537870 133445 538083 133452
rect 536142 133312 536355 133320
rect 536142 133254 536151 133312
rect 536348 133254 536355 133312
rect 536142 133245 536355 133254
rect 534339 133110 534552 133120
rect 534339 133052 534348 133110
rect 534545 133052 534552 133110
rect 534339 133045 534552 133052
rect 534087 132912 534300 132920
rect 534087 132854 534096 132912
rect 534293 132854 534300 132912
rect 534087 132845 534300 132854
rect 533801 132711 534014 132720
rect 533801 132653 533808 132711
rect 534005 132653 534014 132711
rect 533801 132645 534014 132653
rect 533519 132510 533732 132520
rect 533519 132452 533528 132510
rect 533725 132452 533732 132510
rect 533519 132445 533732 132452
rect 533603 132390 533663 132445
rect 533885 132390 533945 132645
rect 534169 132390 534229 132845
rect 534417 132390 534477 133045
rect 536217 132390 536281 133245
rect 537953 132390 538017 133445
rect 551833 132676 551907 134619
rect 551833 132602 583688 132676
rect 533287 132101 583131 132161
rect 452177 112365 452266 113100
rect 456081 112365 456177 113100
rect 452177 89388 456177 112365
rect 583071 94818 583131 132101
rect 583614 96003 583688 132602
rect 584320 96003 585600 96030
rect 583614 95929 583967 96003
rect 584057 95929 585600 96003
rect 584320 95918 585600 95929
rect 584320 94818 585600 94848
rect 583071 94758 585600 94818
rect 584320 94736 585600 94758
rect 584320 93554 584800 93666
rect 584320 92372 584800 92484
rect 452177 88492 452241 89388
rect 456105 88492 456177 89388
rect 290073 30905 290992 30949
rect 290073 30361 290122 30905
rect 290933 30682 290992 30905
rect 290933 30361 290994 30682
rect 290073 30317 290994 30361
rect 7329 22000 285926 22229
rect 3528 18157 4384 18189
rect 3528 17976 3562 18157
rect 1114 17822 3562 17976
rect 0 17710 3562 17822
rect 1114 17563 3562 17710
rect 3528 17264 3562 17563
rect 4344 17264 4384 18157
rect 3528 17233 4384 17264
rect 290074 18165 290994 30317
rect 452177 27991 456177 88492
rect 488832 78206 489758 78234
rect 488832 77954 488864 78206
rect 489714 78188 489758 78206
rect 489714 78174 512103 78188
rect 489714 77972 511606 78174
rect 512088 77972 512103 78174
rect 489714 77954 512103 77972
rect 488832 77922 489758 77954
rect 488770 74217 489966 74243
rect 488770 73965 488810 74217
rect 489925 74186 489966 74217
rect 489925 74171 512094 74186
rect 489925 74031 511558 74171
rect 512077 74031 512094 74171
rect 489925 74016 512094 74031
rect 489925 73965 489966 74016
rect 488770 73936 489966 73965
rect 584320 51344 585600 51372
rect 582433 51277 583665 51344
rect 583752 51277 585600 51344
rect 513831 47212 513909 47227
rect 513831 46976 513838 47212
rect 513899 47042 513909 47212
rect 515337 47220 515415 47235
rect 515337 47042 515344 47220
rect 513899 46984 515344 47042
rect 515405 46984 515415 47220
rect 513899 46978 515415 46984
rect 513899 46976 513909 46978
rect 513831 46966 513909 46976
rect 515337 46974 515415 46978
rect 513521 46308 513621 46321
rect 513521 46055 513539 46308
rect 513603 46055 513621 46308
rect 513521 46036 513621 46055
rect 513546 42037 513613 46036
rect 522986 43472 523046 45871
rect 523666 43731 523726 45866
rect 523584 43723 523815 43731
rect 523584 43664 523599 43723
rect 523806 43664 523815 43723
rect 523584 43655 523815 43664
rect 523666 43627 523726 43655
rect 522986 43452 523335 43472
rect 522986 43386 522999 43452
rect 523317 43386 523335 43452
rect 522986 43370 523335 43386
rect 522986 43365 523046 43370
rect 525026 42277 525086 45903
rect 525706 43931 525766 45861
rect 527066 44131 527126 45866
rect 530853 44331 530913 45857
rect 531203 44531 531263 45857
rect 531511 44731 531571 45857
rect 533590 44931 533654 45861
rect 534187 45131 534247 45857
rect 558669 45554 558783 45925
rect 582433 45554 582509 51277
rect 584320 51260 585600 51277
rect 584320 50160 585600 50190
rect 558669 45481 582509 45554
rect 582620 50091 585600 50160
rect 560829 45366 561153 45372
rect 582620 45366 582689 50091
rect 584320 50078 585600 50091
rect 584320 48896 584800 49008
rect 584320 47714 584800 47826
rect 560829 45357 582689 45366
rect 560829 45301 560845 45357
rect 561136 45301 582689 45357
rect 560829 45297 582689 45301
rect 560829 45289 561153 45297
rect 534085 45124 534316 45131
rect 534085 45065 534097 45124
rect 534304 45065 534316 45124
rect 534085 45055 534316 45065
rect 533496 44922 533727 44931
rect 533496 44863 533511 44922
rect 533718 44863 533727 44922
rect 533496 44855 533727 44863
rect 531414 44723 531645 44731
rect 531414 44664 531429 44723
rect 531636 44664 531645 44723
rect 531414 44655 531645 44664
rect 531111 44523 531342 44531
rect 531111 44464 531124 44523
rect 531331 44464 531342 44523
rect 531111 44455 531342 44464
rect 530758 44323 530989 44331
rect 530758 44264 530771 44323
rect 530978 44264 530989 44323
rect 530758 44255 530989 44264
rect 526976 44123 527207 44131
rect 526976 44064 526989 44123
rect 527196 44064 527207 44123
rect 526976 44055 527207 44064
rect 525615 43923 525846 43931
rect 525615 43864 525627 43923
rect 525834 43864 525846 43923
rect 525615 43855 525846 43864
rect 525706 43627 525766 43855
rect 527066 43627 527126 44055
rect 530853 43627 530913 44255
rect 531203 43627 531263 44455
rect 531511 43627 531571 44655
rect 533590 43627 533654 44855
rect 534187 43627 534247 45055
rect 579433 42523 579551 42545
rect 579433 42277 579450 42523
rect 525026 42203 579450 42277
rect 579433 42199 579450 42203
rect 579522 42199 579551 42523
rect 579433 42173 579551 42199
rect 579104 42037 579222 42048
rect 513546 42026 579223 42037
rect 513546 41963 579123 42026
rect 579104 41702 579123 41963
rect 579195 41963 579223 42026
rect 579195 41702 579222 41963
rect 579104 41676 579222 41702
rect 582047 27991 583234 27996
rect 452177 27953 583249 27991
rect 452177 27654 582111 27953
rect 583186 27654 583249 27953
rect 452177 27602 583249 27654
rect 579118 26872 579240 26894
rect 579118 26514 579140 26872
rect 579213 26514 579240 26872
rect 579118 26494 579240 26514
rect 579421 26871 579543 26897
rect 579421 26513 579438 26871
rect 579511 26513 579543 26871
rect 579421 26497 579543 26513
rect 579750 26872 579872 26898
rect 579750 26514 579770 26872
rect 579843 26514 579872 26872
rect 579750 26498 579872 26514
rect 580115 26872 580237 26897
rect 580115 26514 580133 26872
rect 580206 26514 580237 26872
rect 290074 17259 290103 18165
rect 290967 17259 290994 18165
rect 290074 17234 290994 17259
rect 0 16528 1280 16640
rect 460160 16174 460330 16196
rect 460160 15816 460182 16174
rect 460314 15898 460330 16174
rect 563626 15898 563756 15912
rect 460314 15816 563640 15898
rect 460160 15802 563640 15816
rect 460160 15792 460330 15802
rect 456270 15732 456558 15774
rect 800 15346 1280 15458
rect 181943 14965 182423 14982
rect 181943 14869 181967 14965
rect 182409 14869 182423 14965
rect 456270 14942 456314 15732
rect 456522 15544 456558 15732
rect 456522 15448 563038 15544
rect 563626 15502 563640 15802
rect 563748 15802 563764 15898
rect 563748 15502 563756 15802
rect 563626 15478 563756 15502
rect 456522 14942 456558 15448
rect 562942 15230 563038 15448
rect 562942 15198 564046 15230
rect 562942 15134 563932 15198
rect 456270 14892 456558 14942
rect 181943 14855 182423 14869
rect 800 14164 1280 14276
rect 0 12982 1280 13094
rect 0 11800 1280 11912
rect 800 10618 1280 10730
rect 800 9436 1280 9548
rect 0 8254 1280 8366
rect 182149 7460 182247 14855
rect 563906 14808 563932 15134
rect 564020 14808 564046 15198
rect 563906 14778 564046 14808
rect 280227 11091 280448 11093
rect 288826 11091 289047 11093
rect 260952 11088 289047 11091
rect 260952 11032 280236 11088
rect 280439 11032 288835 11088
rect 289038 11032 289047 11088
rect 260952 11027 289047 11032
rect 279879 10963 280100 10965
rect 288452 10963 288673 10965
rect 260952 10960 288997 10963
rect 260952 10904 279888 10960
rect 280091 10904 288461 10960
rect 288664 10904 288997 10960
rect 260952 10899 288997 10904
rect 279510 10835 279731 10837
rect 288248 10835 288469 10837
rect 260952 10832 288997 10835
rect 260952 10776 279573 10832
rect 279722 10776 288257 10832
rect 288460 10776 288997 10832
rect 260952 10771 288997 10776
rect 279186 10707 279407 10709
rect 288053 10707 288274 10709
rect 260952 10704 288997 10707
rect 260952 10648 279262 10704
rect 279398 10648 288062 10704
rect 288265 10648 288997 10704
rect 260952 10643 288997 10648
rect 298868 10678 299194 10694
rect 298868 10620 298896 10678
rect 299168 10670 299194 10678
rect 569644 10676 569964 10692
rect 569644 10670 569672 10676
rect 299168 10620 569672 10670
rect 298868 10600 569672 10620
rect 569644 10590 569672 10600
rect 569944 10590 569964 10676
rect 278837 10579 279058 10582
rect 287856 10579 288077 10581
rect 260952 10577 288997 10579
rect 260952 10521 278859 10577
rect 279049 10576 288997 10577
rect 279049 10521 287865 10576
rect 260952 10520 287865 10521
rect 288068 10520 288997 10576
rect 569644 10574 569964 10590
rect 297350 10532 297571 10535
rect 403147 10532 403368 10535
rect 260952 10515 288997 10520
rect 297282 10530 424679 10532
rect 297282 10474 297359 10530
rect 297562 10474 403156 10530
rect 403359 10474 424679 10530
rect 297282 10468 424679 10474
rect 278479 10451 278700 10452
rect 287654 10451 287875 10453
rect 260952 10448 288997 10451
rect 260952 10447 287663 10448
rect 260952 10391 278570 10447
rect 278691 10392 287663 10447
rect 287866 10392 288997 10448
rect 297546 10404 297767 10407
rect 406701 10404 406922 10407
rect 278691 10391 288997 10392
rect 260952 10387 288997 10391
rect 297282 10402 424679 10404
rect 278479 10386 278700 10387
rect 297282 10346 297555 10402
rect 297758 10346 406710 10402
rect 406913 10346 424679 10402
rect 297282 10340 424679 10346
rect 278145 10323 278366 10324
rect 287455 10323 287676 10325
rect 260952 10320 288997 10323
rect 260952 10319 287464 10320
rect 260952 10263 278154 10319
rect 278357 10264 287464 10319
rect 287667 10264 288997 10320
rect 297744 10276 297965 10279
rect 410259 10276 410480 10279
rect 278357 10263 288997 10264
rect 260952 10259 288997 10263
rect 297282 10274 424679 10276
rect 278145 10258 278366 10259
rect 297282 10218 297753 10274
rect 297956 10218 410268 10274
rect 410471 10218 424679 10274
rect 297282 10212 424679 10218
rect 275208 10195 275429 10196
rect 287246 10195 287467 10198
rect 260952 10193 288997 10195
rect 260952 10191 287255 10193
rect 260952 10135 275217 10191
rect 275420 10137 287255 10191
rect 287458 10137 288997 10193
rect 297951 10148 298172 10150
rect 413807 10148 414028 10149
rect 275420 10135 288997 10137
rect 260952 10131 288997 10135
rect 297282 10145 424679 10148
rect 275208 10130 275429 10131
rect 297282 10089 297960 10145
rect 298163 10144 424679 10145
rect 298163 10089 413816 10144
rect 297282 10088 413816 10089
rect 414019 10088 424679 10144
rect 297282 10084 424679 10088
rect 413807 10083 414028 10084
rect 271654 10067 271878 10070
rect 287060 10067 287281 10069
rect 260952 10065 288997 10067
rect 260952 10009 271663 10065
rect 271866 10064 288997 10065
rect 271866 10009 287069 10064
rect 260952 10008 287069 10009
rect 287272 10008 288997 10064
rect 298149 10020 298370 10023
rect 417344 10020 417565 10022
rect 260952 10003 288997 10008
rect 297282 10018 424679 10020
rect 297282 9962 298158 10018
rect 298361 10017 424679 10018
rect 298361 9962 417353 10017
rect 297282 9961 417353 9962
rect 417556 9961 424679 10017
rect 297282 9956 424679 9961
rect 268130 9939 268351 9942
rect 286857 9939 287078 9941
rect 260952 9937 288997 9939
rect 260952 9881 268139 9937
rect 268342 9936 288997 9937
rect 268342 9881 286866 9936
rect 260952 9880 286866 9881
rect 287069 9880 288997 9936
rect 298345 9892 298566 9895
rect 420880 9892 421101 9893
rect 260952 9875 288997 9880
rect 297282 9890 424679 9892
rect 297282 9834 298354 9890
rect 298557 9888 424679 9890
rect 298557 9834 420889 9888
rect 297282 9832 420889 9834
rect 421092 9832 424679 9888
rect 297282 9828 424679 9832
rect 420880 9827 421101 9828
rect 264553 9811 264774 9812
rect 286670 9811 286891 9813
rect 260952 9808 288997 9811
rect 260952 9807 286679 9808
rect 260952 9751 264562 9807
rect 264765 9752 286679 9807
rect 286882 9752 288997 9808
rect 298541 9764 298762 9767
rect 424454 9764 424675 9766
rect 264765 9751 288997 9752
rect 260952 9747 288997 9751
rect 297282 9762 424679 9764
rect 264553 9746 264774 9747
rect 297282 9706 298550 9762
rect 298753 9761 424679 9762
rect 298753 9706 424463 9761
rect 297282 9705 424463 9706
rect 424666 9705 424679 9761
rect 297282 9700 424679 9705
rect 261008 9683 261229 9685
rect 286452 9683 286673 9685
rect 260952 9680 288997 9683
rect 260952 9624 261017 9680
rect 261220 9624 286461 9680
rect 286664 9624 288997 9680
rect 260952 9619 288997 9624
rect 181525 7436 182295 7460
rect 181525 7340 181554 7436
rect 182266 7340 182295 7436
rect 181525 7316 182295 7340
rect 0 7072 1280 7184
rect 800 5890 1280 6002
rect 800 4708 1280 4820
rect 579155 4797 579222 26494
rect 579448 9530 579515 26497
rect 579777 14241 579838 26498
rect 580115 26497 580237 26514
rect 580420 26879 580542 26900
rect 580420 26521 580440 26879
rect 580513 26521 580542 26879
rect 580420 26500 580542 26521
rect 580137 18981 580198 26497
rect 580456 23705 580517 26500
rect 582966 25125 583171 25153
rect 582966 24613 583000 25125
rect 583140 24878 583171 25125
rect 584320 24878 585600 24914
rect 583140 24817 583804 24878
rect 583889 24817 585600 24878
rect 583140 24613 583171 24817
rect 584320 24802 585600 24817
rect 582966 24581 583171 24613
rect 584320 23705 585600 23732
rect 580452 23644 585600 23705
rect 584320 23620 585600 23644
rect 584320 22438 584800 22550
rect 584320 21256 584800 21368
rect 582960 20364 583165 20403
rect 582960 19852 582991 20364
rect 583131 20142 583165 20364
rect 584320 20142 585600 20186
rect 583131 20081 583801 20142
rect 583886 20081 585600 20142
rect 583131 19852 583165 20081
rect 584320 20074 585600 20081
rect 582960 19831 583165 19852
rect 584320 18981 585600 19004
rect 580137 18920 585600 18981
rect 584320 18892 585600 18920
rect 584320 17710 584800 17822
rect 584320 16528 584800 16640
rect 582966 15647 583171 15678
rect 582966 15135 583004 15647
rect 583144 15416 583171 15647
rect 584320 15416 585600 15458
rect 583144 15355 583847 15416
rect 583932 15355 585600 15416
rect 583144 15135 583171 15355
rect 584320 15346 585600 15355
rect 582966 15106 583171 15135
rect 584320 14241 585600 14276
rect 579777 14180 585600 14241
rect 584320 14164 585600 14180
rect 584320 12982 584800 13094
rect 584320 11800 584800 11912
rect 582976 10933 583181 10963
rect 582976 10421 583002 10933
rect 583142 10716 583181 10933
rect 584320 10716 585600 10730
rect 583142 10635 583803 10716
rect 583891 10635 585600 10716
rect 583142 10421 583181 10635
rect 584320 10618 585600 10635
rect 582976 10391 583181 10421
rect 584320 9530 585600 9548
rect 579448 9463 585600 9530
rect 584320 9436 585600 9463
rect 584320 8254 584800 8366
rect 584320 7072 584800 7184
rect 582970 6190 583175 6213
rect 582970 5664 583003 6190
rect 583137 5977 583175 6190
rect 584320 5977 585600 6002
rect 583137 5896 583839 5977
rect 583927 5896 585600 5977
rect 583137 5664 583175 5896
rect 584320 5890 585600 5896
rect 582970 5641 583175 5664
rect 584320 4797 585600 4820
rect 579155 4730 585600 4797
rect 584320 4708 585600 4730
rect 0 3526 1280 3638
rect 584320 3526 584800 3638
rect 0 2344 1280 2456
rect 584320 2344 584800 2456
<< rmetal3 >>
rect 1288 376754 1353 376866
rect 1444 33126 1626 33416
rect 583582 590272 583722 590384
rect 583574 500850 583714 500962
rect 583522 320362 583662 320474
rect 583756 275940 583896 276052
rect 583967 95929 584057 96003
rect 583665 51277 583752 51344
rect 583804 24817 583889 24878
rect 583801 20081 583886 20142
rect 583847 15355 583932 15416
rect 583803 10635 583891 10716
rect 583839 5896 583927 5977
<< via3 >>
rect 3472 644833 8318 649314
rect 3494 634779 8340 639260
rect 4054 560414 9132 564868
rect 4066 550426 9144 554880
rect 100018 504650 102298 507328
rect 28395 486659 38334 492430
rect 18241 478121 18645 479537
rect 6256 470365 12269 475393
rect 7523 461352 8290 461984
rect 5436 455115 6072 456528
rect 43381 443121 44947 452040
rect 104310 446394 106146 448182
rect 6378 429877 7086 430832
rect 11697 427828 13585 428240
rect 8126 384475 9182 384757
rect 73831 384033 74622 384777
rect 8553 382858 9115 383290
rect 8241 381897 9368 382289
rect 7617 379740 9223 379992
rect 7609 378984 9228 379239
rect 1392 376729 2159 376882
rect 59828 363848 60326 364712
rect 116072 345626 118072 347766
rect 4983 339220 5982 339653
rect 11146 335652 11723 336581
rect 6789 334800 7923 335356
rect 3091 311780 3736 314581
rect 25702 318190 26022 318928
rect 7588 306618 7747 307000
rect 50036 310072 50460 310650
rect 10019 307782 10174 308203
rect 10018 302398 10174 302786
rect 10668 305956 10827 306338
rect 50036 306142 50462 306986
rect 5290 296044 6335 296534
rect 8908 292471 9750 293051
rect 7102 291597 8352 292119
rect 11839 302797 12083 302878
rect 11835 302596 12079 302677
rect 9820 287428 10389 287991
rect 5242 286612 6400 287221
rect 128918 652362 132733 653097
rect 136910 653988 140725 654723
rect 136986 639691 140674 644370
rect 129074 589599 132598 595069
rect 128910 562358 132725 563093
rect 128924 472150 132768 475246
rect 128923 382381 132755 383136
rect 128918 379827 132762 380144
rect 128962 376582 132722 377026
rect 128893 363838 132628 364692
rect 128934 310102 132738 310649
rect 128935 292378 132733 293105
rect 7809 285650 8396 286306
rect 122182 284192 124562 286830
rect 4310 215890 9440 220396
rect 10348 218145 11403 220037
rect 4284 205852 9414 210358
rect 128929 202363 132761 203118
rect 3756 173829 8602 178310
rect 129023 168834 132621 173511
rect 3676 163839 8522 168320
rect 122080 116572 124173 117189
rect 8320 109813 10127 113162
rect 128914 112351 132746 113106
rect 4550 104052 6568 107789
rect 7550 84414 9045 85317
rect 9045 84414 9901 85317
rect 9901 84414 11060 85317
rect 5768 82240 9278 83143
rect 128916 84353 132725 85335
rect 3917 78534 4887 79506
rect 128967 53284 132708 56959
rect 5712 38923 6434 39422
rect 113278 31500 118898 32468
rect 136911 563973 140726 564708
rect 136918 476568 140733 477303
rect 137099 391475 140611 401010
rect 136941 383956 140773 384711
rect 136999 378850 140729 379269
rect 136912 361328 140668 362468
rect 136918 309106 140746 309624
rect 136946 293979 140744 294706
rect 136923 203968 140755 204723
rect 146008 143960 148318 146268
rect 136938 113982 140770 114737
rect 136942 82204 140751 83186
rect 511510 693868 516020 698944
rect 521554 693856 526064 698932
rect 263662 653984 265591 654713
rect 321200 653975 323129 654704
rect 245788 652377 247717 653106
rect 339074 652368 341003 653097
rect 422844 604042 425668 606998
rect 283246 567566 284368 567908
rect 263662 563984 265591 564713
rect 245788 562377 247717 563106
rect 263662 476584 265591 477313
rect 245788 472377 247717 473106
rect 263662 383984 265591 384713
rect 245788 382377 247717 383106
rect 321200 563975 323129 564704
rect 339074 562368 341003 563097
rect 284414 477428 284791 478603
rect 263662 293984 265591 294713
rect 245788 292377 247717 293106
rect 283572 293605 283964 295162
rect 321200 473975 323129 474704
rect 339074 472368 341003 473097
rect 286018 385768 287145 386083
rect 321200 383975 323129 384704
rect 339074 382368 341003 383097
rect 339074 294368 341003 295097
rect 321212 292187 323141 292916
rect 423834 497872 424381 499533
rect 426592 428204 428498 430286
rect 421370 292005 422855 292454
rect 423897 291416 425382 291865
rect 289130 288524 290210 288789
rect 289114 287037 290194 287302
rect 289110 286396 290190 286661
rect 299365 285048 299882 285969
rect 300312 285038 300829 285959
rect 284796 278144 285034 278775
rect 285179 276044 285438 276685
rect 285676 273948 285943 274532
rect 427136 284006 430734 287604
rect 444265 653958 448080 654693
rect 444374 635697 448011 640383
rect 444283 563978 448098 564713
rect 438977 386616 439074 386918
rect 452277 652358 456092 653093
rect 573828 640732 578952 645170
rect 573842 630762 578966 635200
rect 508882 594750 510528 595050
rect 513911 593259 520276 609778
rect 510907 570179 518330 576926
rect 452281 562359 456096 563094
rect 452220 500838 456132 500973
rect 452284 491981 456101 492374
rect 444298 491240 448085 491676
rect 444287 473967 448102 474702
rect 444261 383975 448076 384710
rect 444363 355510 448074 356155
rect 440123 354020 440396 355012
rect 444353 309389 448020 310336
rect 444258 297698 448110 298616
rect 444240 295951 448055 296686
rect 442709 276714 442977 277307
rect 440930 273577 441236 274403
rect 433885 209657 434271 211499
rect 436894 209632 437280 211474
rect 164278 205964 165881 206339
rect 263662 203984 265591 204713
rect 245788 202377 247717 203106
rect 321200 203975 323129 204704
rect 423193 205481 424985 205978
rect 433860 204374 434276 206427
rect 436868 204358 437284 206411
rect 339074 202368 341003 203097
rect 423476 195753 424871 196209
rect 164579 116604 166211 117154
rect 431353 163637 434495 167041
rect 263662 113984 265591 114713
rect 245788 112377 247717 113106
rect 159964 63802 162104 66158
rect 321200 113975 323129 114704
rect 339074 112368 341003 113097
rect 440954 155284 441137 156125
rect 442705 156171 442983 156796
rect 444285 201720 448100 202455
rect 444303 179958 448071 180774
rect 452283 472385 456098 473120
rect 573573 585613 574366 586727
rect 577145 583409 577661 584173
rect 575644 551600 580768 556038
rect 575630 541566 580754 546004
rect 460928 500842 461800 500977
rect 576075 496743 576616 498421
rect 575013 495447 575808 496291
rect 576790 493993 577757 494849
rect 578317 492070 579412 492276
rect 578266 491321 579420 491568
rect 476138 425383 479384 434151
rect 466355 410038 473541 412620
rect 580603 384268 581287 384575
rect 452289 382392 456104 383127
rect 582944 365988 583273 368196
rect 580208 360563 581211 361187
rect 452253 357386 456061 358012
rect 575167 357360 576400 358018
rect 575129 355501 576287 356137
rect 579107 354393 580386 354648
rect 567177 315844 568123 316809
rect 569330 314111 569965 315568
rect 571103 313895 572537 314309
rect 452287 306064 456063 306969
rect 565640 309073 566219 310201
rect 564258 305360 564610 306470
rect 581414 297785 581521 298423
rect 582339 297784 582446 298422
rect 513273 295445 513751 295774
rect 452291 294384 456106 295119
rect 452238 292590 456120 293534
rect 495054 283618 495406 283932
rect 497633 279505 498017 279858
rect 567218 271604 568058 272396
rect 578316 270535 579119 270783
rect 578330 269456 579103 269758
rect 564172 267178 564723 267662
rect 565565 265643 566309 266037
rect 525018 250571 525156 250793
rect 525018 249837 525156 250059
rect 529560 250354 529698 250576
rect 529935 250338 530073 250560
rect 530303 250362 530441 250584
rect 529549 249566 529687 249788
rect 529940 249573 530078 249795
rect 530288 249586 530426 249808
rect 574934 236252 580058 240690
rect 574962 226222 580086 230660
rect 452266 199609 456081 200344
rect 574896 192412 580020 196850
rect 452333 187251 455990 191899
rect 574908 182368 580032 186806
rect 452276 176624 456058 177478
rect 444260 113976 448075 114711
rect 444290 91356 448055 92247
rect 442690 77894 443023 78912
rect 440192 73811 440394 74403
rect 436136 63691 439734 67289
rect 137083 31547 140503 40865
rect 129020 23480 132614 28804
rect 492662 156162 493194 156342
rect 494004 155582 494639 155736
rect 575156 147818 580280 152256
rect 575102 137756 580226 142194
rect 452266 112365 456081 113100
rect 452241 88492 456105 89388
rect 3562 17264 4344 18157
rect 488864 77954 489714 78206
rect 488810 73965 489925 74217
rect 290103 17259 290967 18165
<< metal4 >>
rect 166394 703100 171394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 330094 703100 335094 704800
rect 511354 698944 526180 699076
rect 511354 693868 511510 698944
rect 516020 698932 526180 698944
rect 516020 693868 516456 698932
rect 511354 693856 516456 693868
rect 520966 693856 521554 698932
rect 526064 693856 526180 698932
rect 511354 693672 526180 693856
rect 263426 654796 265741 654863
rect 128043 654723 265741 654796
rect 128043 653988 136910 654723
rect 140725 654713 265741 654723
rect 140725 653988 263662 654713
rect 128043 653984 263662 653988
rect 265591 653984 265741 654713
rect 128043 653892 265741 653984
rect 263426 653791 265741 653892
rect 321050 654787 323365 654854
rect 321050 654704 456383 654787
rect 321050 653975 321200 654704
rect 323129 654693 456383 654704
rect 323129 653975 444265 654693
rect 321050 653958 444265 653975
rect 448080 653958 456383 654693
rect 321050 653883 456383 653958
rect 321050 653782 323365 653883
rect 245574 653196 247889 653256
rect 128043 653106 247904 653196
rect 338902 653187 341217 653247
rect 128043 653097 245788 653106
rect 128043 652362 128918 653097
rect 132733 652377 245788 653097
rect 247717 652377 247904 653106
rect 132733 652362 247904 652377
rect 128043 652292 247904 652362
rect 338887 653097 456383 653187
rect 338887 652368 339074 653097
rect 341003 653093 456383 653097
rect 341003 652368 452277 653093
rect 338887 652358 452277 652368
rect 456092 652358 456383 653093
rect 245574 652184 247889 652292
rect 338887 652283 456383 652358
rect 338902 652175 341217 652283
rect 3308 649314 8544 649486
rect 3308 644833 3472 649314
rect 8318 644833 8544 649314
rect 3308 644534 8544 644833
rect 573700 645170 579138 645386
rect 3308 644370 141468 644534
rect 3308 639691 136986 644370
rect 140674 639691 141468 644370
rect 573700 640732 573828 645170
rect 578952 640732 579138 645170
rect 573700 640538 579138 640732
rect 3308 639534 141468 639691
rect 443754 640383 579138 640538
rect 3308 639260 8544 639534
rect 3308 634779 3494 639260
rect 8340 634779 8544 639260
rect 443754 635697 444374 640383
rect 448011 635697 579138 640383
rect 443754 635538 579138 635697
rect 3308 634618 8544 634779
rect 573700 635200 579138 635538
rect 573700 630762 573842 635200
rect 578966 630762 579138 635200
rect 573700 630566 579138 630762
rect 98259 601186 169654 610368
rect 417050 610315 515494 610324
rect 417050 609778 520733 610315
rect 417050 606998 513911 609778
rect 417050 604042 422844 606998
rect 425668 604042 513911 606998
rect 417050 601142 513911 604042
rect 128823 595069 132844 595370
rect 128823 594559 129074 595069
rect 98259 593599 129074 594559
rect 128823 589599 129074 593599
rect 132598 589599 132844 595069
rect 508780 595050 510602 595116
rect 513415 595070 513911 601142
rect 508780 595028 508882 595050
rect 128823 589258 132844 589599
rect 422781 594750 508882 595028
rect 510528 594750 510602 595050
rect 422781 594726 510602 594750
rect 513414 594741 513911 595070
rect 283206 567908 284412 567940
rect 283206 567566 283246 567908
rect 284368 567895 284412 567908
rect 422781 567895 423083 594726
rect 508780 594670 510602 594726
rect 513415 593259 513911 594741
rect 520276 593259 520733 609778
rect 513415 592789 520733 593259
rect 573463 586727 574467 586813
rect 573463 585613 573573 586727
rect 574366 585613 574467 586727
rect 573463 585534 574467 585613
rect 466103 577278 518844 577547
rect 466103 569837 466468 577278
rect 473449 576926 518844 577278
rect 473449 570179 510907 576926
rect 518330 570179 518844 576926
rect 473449 569837 518844 570179
rect 466103 569612 518844 569837
rect 284368 567593 423083 567895
rect 284368 567566 284412 567593
rect 283206 567534 284412 567566
rect 3906 564868 9344 565044
rect 3906 560414 4054 564868
rect 9132 560414 9344 564868
rect 263426 564796 265741 564863
rect 127952 564713 265741 564796
rect 127952 564708 263662 564713
rect 127952 563973 136911 564708
rect 140726 563984 263662 564708
rect 265591 563984 265741 564713
rect 140726 563973 265741 563984
rect 127952 563892 265741 563973
rect 263426 563791 265741 563892
rect 321050 564787 323365 564854
rect 321050 564713 456394 564787
rect 321050 564704 444283 564713
rect 321050 563975 321200 564704
rect 323129 563978 444283 564704
rect 448098 563978 456394 564713
rect 323129 563975 456394 563978
rect 321050 563883 456394 563975
rect 321050 563782 323365 563883
rect 245574 563196 247889 563256
rect 127952 563106 247904 563196
rect 338902 563187 341217 563247
rect 127952 563093 245788 563106
rect 127952 562358 128910 563093
rect 132725 562377 245788 563093
rect 247717 562377 247904 563106
rect 132725 562358 247904 562377
rect 127952 562292 247904 562358
rect 338887 563097 456394 563187
rect 338887 562368 339074 563097
rect 341003 563094 456394 563097
rect 341003 562368 452281 563094
rect 338887 562359 452281 562368
rect 456096 562359 456394 563094
rect 245574 562184 247889 562292
rect 338887 562283 456394 562359
rect 338902 562175 341217 562283
rect 3906 560048 9344 560414
rect 3906 555362 4066 560048
rect 9170 555362 9344 560048
rect 3906 554880 9344 555362
rect 3906 550426 4066 554880
rect 9144 550426 9344 554880
rect 3906 550224 9344 550426
rect 466125 560021 473749 560331
rect 466125 553646 466599 560021
rect 473439 553646 473749 560021
rect 466125 530621 473749 553646
rect 466125 523885 466547 530621
rect 473413 523885 473749 530621
rect 573472 530016 574169 585534
rect 577090 584230 577539 584238
rect 577087 584173 577726 584230
rect 577087 583409 577145 584173
rect 577661 583409 577726 584173
rect 577087 583360 577726 583409
rect 577090 556170 577539 583360
rect 575502 556038 580940 556170
rect 575502 551600 575644 556038
rect 580768 551600 580940 556038
rect 575502 550970 580940 551600
rect 575502 546532 575622 550970
rect 580746 546532 580940 550970
rect 575502 546004 580940 546532
rect 575502 541566 575630 546004
rect 580754 541566 580940 546004
rect 575502 541350 580940 541566
rect 572142 529912 574258 530016
rect 572142 527565 572241 529912
rect 574152 527565 574258 529912
rect 572142 527489 574258 527565
rect 466125 523522 473749 523885
rect 60811 507328 169654 510368
rect 60811 504650 100018 507328
rect 102298 504650 169654 507328
rect 417050 505142 486115 514324
rect 60811 501186 169654 504650
rect 573472 502532 574169 527489
rect 573472 501835 576687 502532
rect 60811 494403 69993 501186
rect 452180 500977 461847 501013
rect 452180 500973 460928 500977
rect 452180 500838 452220 500973
rect 456132 500842 460928 500973
rect 461800 500842 461847 500977
rect 456132 500838 461847 500842
rect 452180 500810 461847 500838
rect 423770 499533 424448 499585
rect 423770 497872 423834 499533
rect 424381 498942 424448 499533
rect 424381 498488 575615 498942
rect 424381 497872 424448 498488
rect 423770 497813 424448 497872
rect 575161 496393 575615 498488
rect 575990 498421 576687 501835
rect 575990 496743 576075 498421
rect 576616 496743 576687 498421
rect 575990 496650 576687 496743
rect 574914 496291 575907 496393
rect 574914 495447 575013 496291
rect 575808 495447 575907 496291
rect 574914 495358 575907 495447
rect 575161 495356 575615 495358
rect 577090 494922 577539 541350
rect 27578 492430 69993 494403
rect 576700 494849 577862 494922
rect 576700 493993 576790 494849
rect 577757 493993 577862 494849
rect 576700 493929 577862 493993
rect 27578 486659 28395 492430
rect 38334 486659 69993 492430
rect 452154 492374 456203 492443
rect 452154 491981 452284 492374
rect 456101 492320 456203 492374
rect 456101 492276 579461 492320
rect 456101 492070 578317 492276
rect 579412 492070 579461 492276
rect 456101 492034 579461 492070
rect 456101 491981 456203 492034
rect 578266 492032 579461 492034
rect 452154 491916 456203 491981
rect 444107 491676 448181 491793
rect 444107 491240 444298 491676
rect 448085 491586 448181 491676
rect 578225 491586 579451 491594
rect 448085 491568 579451 491586
rect 448085 491321 578266 491568
rect 579420 491321 579451 491568
rect 448085 491300 579451 491321
rect 448085 491240 448181 491300
rect 578225 491282 579451 491300
rect 444107 491144 448181 491240
rect 27578 485221 69993 486659
rect 18196 479537 18710 479594
rect 18196 478121 18241 479537
rect 18645 478497 18710 479537
rect 284377 478603 284838 478643
rect 284377 478497 284414 478603
rect 18645 478121 284414 478497
rect 18196 478067 284414 478121
rect 18196 478064 18710 478067
rect 263426 477396 265741 477463
rect 128446 477313 265741 477396
rect 284377 477428 284414 478067
rect 284791 477428 284838 478603
rect 284377 477375 284838 477428
rect 128446 477303 263662 477313
rect 128446 476568 136918 477303
rect 140733 476584 263662 477303
rect 265591 476584 265741 477313
rect 140733 476568 265741 476584
rect 128446 476492 265741 476568
rect 263426 476391 265741 476492
rect 4420 475393 114425 475493
rect 4420 470365 6256 475393
rect 12269 475380 114425 475393
rect 12269 470365 106611 475380
rect 4420 470309 106611 470365
rect 113894 470309 114425 475380
rect 128686 475246 280750 475394
rect 128686 472150 128924 475246
rect 132768 475224 280750 475246
rect 132768 473106 273494 475224
rect 132768 472377 245788 473106
rect 247717 472377 273494 473106
rect 132768 472164 273494 472377
rect 280502 472164 280750 475224
rect 321050 474787 323365 474854
rect 321050 474704 456315 474787
rect 321050 473975 321200 474704
rect 323129 474702 456315 474704
rect 323129 473975 444287 474702
rect 321050 473967 444287 473975
rect 448102 473967 456315 474702
rect 321050 473883 456315 473967
rect 321050 473782 323365 473883
rect 338902 473187 341217 473247
rect 338887 473120 456315 473187
rect 338887 473097 452283 473120
rect 338887 472368 339074 473097
rect 341003 472385 452283 473097
rect 456098 472385 456315 473120
rect 341003 472368 456315 472385
rect 338887 472283 456315 472368
rect 338902 472175 341217 472283
rect 132768 472150 280750 472164
rect 128686 471952 280750 472150
rect 4420 470219 114425 470309
rect 150797 462824 158032 462940
rect 150797 462028 150899 462824
rect 7466 461984 150899 462028
rect 7466 461352 7523 461984
rect 8290 461395 150899 461984
rect 157916 462028 158032 462824
rect 157916 461395 158180 462028
rect 8290 461352 158180 461395
rect 7466 461302 158180 461352
rect 150797 461301 158032 461302
rect 5343 456528 6129 456631
rect 5343 455115 5436 456528
rect 6072 455757 6129 456528
rect 106510 455757 114021 455761
rect 6072 455661 114021 455757
rect 6072 455115 106619 455661
rect 5343 455031 106619 455115
rect 106510 454319 106619 455031
rect 113903 454319 114021 455661
rect 106510 454196 114021 454319
rect 42751 452040 169654 452168
rect 42751 443121 43381 452040
rect 44947 448182 169654 452040
rect 44947 446394 104310 448182
rect 106146 446394 169654 448182
rect 44947 443121 169654 446394
rect 42751 442986 169654 443121
rect 106528 441575 114020 441685
rect 106528 440841 106630 441575
rect 81054 440408 106630 440841
rect 113902 440841 114020 441575
rect 113902 440408 114120 440841
rect 81054 440326 114120 440408
rect 150780 440395 158029 440524
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 6302 429814 7162 429877
rect 6469 427411 7004 429814
rect 81054 428297 81569 440326
rect 106528 440321 114020 440326
rect 150780 439439 150941 440395
rect 11637 428240 81569 428297
rect 11637 427828 11697 428240
rect 13585 427828 81569 428240
rect 11637 427782 81569 427828
rect 82329 439040 150941 439439
rect 157881 439040 158029 440395
rect 82329 438906 158029 439040
rect 82329 438904 157979 438906
rect 82329 427411 82864 438904
rect 6469 426876 82864 427411
rect 417050 434151 479733 434324
rect 417050 430286 476138 434151
rect 417050 428204 426592 430286
rect 428498 428204 476138 430286
rect 417050 425383 476138 428204
rect 479384 425383 479733 434151
rect 417050 425142 479733 425383
rect 466206 412620 473703 412769
rect 466206 410038 466355 412620
rect 473541 410038 473703 412620
rect 466206 409865 473703 410038
rect 136611 401010 167867 401173
rect 136611 391475 137099 401010
rect 140611 400684 167867 401010
rect 140611 391614 163821 400684
rect 167356 391614 167867 400684
rect 140611 391475 167867 391614
rect 136611 391172 167867 391475
rect 106531 387634 114007 387717
rect 106531 387504 106648 387634
rect 68878 387152 106648 387504
rect 68878 384793 69230 387152
rect 106531 387014 106648 387152
rect 113913 387014 114007 387634
rect 106531 386917 114007 387014
rect 438962 386919 439091 386935
rect 120639 386918 482545 386919
rect 120639 386616 438977 386918
rect 439074 386616 482545 386918
rect 120639 386612 482545 386616
rect 8087 384757 69230 384793
rect 8087 384475 8126 384757
rect 9182 384475 69230 384757
rect 8087 384441 69230 384475
rect 73769 384777 74673 384820
rect 73769 384033 73831 384777
rect 74622 384569 74673 384777
rect 120639 384569 120946 386612
rect 438962 386597 439091 386612
rect 285962 386083 287206 386139
rect 285962 386006 286018 386083
rect 74622 384262 120946 384569
rect 124682 385807 286018 386006
rect 74622 384033 74673 384262
rect 73769 383978 74673 384033
rect 8490 383290 9178 383354
rect 8490 382858 8553 383290
rect 9115 383006 9178 383290
rect 124682 383006 124881 385807
rect 285962 385768 286018 385807
rect 287145 385768 287206 386083
rect 285962 385713 287206 385768
rect 263426 384796 265741 384863
rect 128580 384713 265741 384796
rect 128580 384711 263662 384713
rect 128580 383956 136941 384711
rect 140773 383984 263662 384711
rect 265591 383984 265741 384713
rect 321050 384787 323365 384854
rect 321050 384710 456385 384787
rect 321050 384704 444261 384710
rect 321050 384569 321200 384704
rect 321049 384262 321200 384569
rect 140773 383956 265741 383984
rect 128580 383892 265741 383956
rect 263426 383791 265741 383892
rect 321050 383975 321200 384262
rect 323129 383975 444261 384704
rect 448076 383975 456385 384710
rect 482238 384569 482545 386612
rect 580563 384575 581315 384602
rect 580563 384569 580603 384575
rect 482238 384268 580603 384569
rect 581287 384268 581315 384575
rect 482238 384262 581315 384268
rect 580563 384240 581315 384262
rect 321050 383883 456385 383975
rect 321050 383782 323365 383883
rect 245574 383196 247889 383256
rect 9115 382858 124881 383006
rect 8490 382807 124881 382858
rect 128580 383136 247904 383196
rect 338902 383187 341217 383247
rect 128580 382381 128923 383136
rect 132755 383106 247904 383136
rect 132755 382381 245788 383106
rect 128580 382377 245788 382381
rect 247717 382377 247904 383106
rect 8167 382289 125973 382347
rect 128580 382292 247904 382377
rect 338887 383127 456385 383187
rect 338887 383097 452289 383127
rect 338887 382368 339074 383097
rect 341003 382392 452289 383097
rect 456104 382392 456385 383127
rect 341003 382368 456385 382392
rect 8167 381897 8241 382289
rect 9368 381897 125973 382289
rect 245574 382184 247889 382292
rect 338887 382283 456385 382368
rect 338902 382175 341217 382283
rect 8167 381846 125973 381897
rect 125472 381147 125973 381846
rect 150787 381147 158044 381204
rect 125472 381083 158044 381147
rect 125472 380646 150869 381083
rect 128817 380144 132851 380208
rect 128817 380019 128918 380144
rect 7571 379992 128918 380019
rect 7571 379740 7617 379992
rect 9223 379827 128918 379992
rect 132762 380019 132851 380144
rect 150787 380153 150869 380646
rect 157943 380153 158044 381083
rect 150787 380065 158044 380153
rect 132762 379827 132854 380019
rect 9223 379740 132854 379827
rect 7571 379709 132854 379740
rect 136847 379269 140818 379383
rect 136847 379263 136999 379269
rect 7566 379239 136999 379263
rect 7566 378984 7609 379239
rect 9228 378984 136999 379239
rect 7566 378955 136999 378984
rect 136847 378850 136999 378955
rect 140729 379263 140818 379269
rect 140729 378955 140845 379263
rect 140729 378850 140818 378955
rect 136847 378723 140818 378850
rect 128879 377026 132795 377076
rect 128879 376909 128962 377026
rect 1363 376882 128962 376909
rect 1363 376729 1392 376882
rect 2159 376729 128962 376882
rect 1363 376706 128962 376729
rect 128879 376582 128962 376706
rect 132722 376582 132795 377026
rect 128879 376525 132795 376582
rect 417050 371142 485757 380324
rect 4935 369733 158189 369749
rect 4842 369602 158189 369733
rect 4842 366820 150962 369602
rect 157821 366820 158189 369602
rect 466227 368377 473688 368506
rect 466227 367103 466376 368377
rect 473507 368077 473688 368377
rect 582908 368196 583306 368262
rect 582908 368077 582944 368196
rect 473507 367329 582944 368077
rect 473507 367103 473688 367329
rect 466227 366922 473688 367103
rect 4842 366667 158189 366820
rect 4842 339653 6115 366667
rect 582908 365988 582944 367329
rect 583273 365988 583306 368196
rect 582908 365946 583306 365988
rect 4842 339220 4983 339653
rect 5982 339220 6115 339653
rect 4842 332034 6115 339220
rect 10039 364712 132687 364758
rect 10039 363848 59828 364712
rect 60326 364692 132687 364712
rect 60326 363848 128893 364692
rect 10039 363838 128893 363848
rect 132628 363838 132687 364692
rect 10039 363790 132687 363838
rect 6704 335356 8008 335437
rect 6704 334800 6789 335356
rect 7923 335271 8008 335356
rect 10039 335271 10526 363790
rect 11113 362468 140772 362536
rect 11113 361328 136912 362468
rect 140668 361328 140772 362468
rect 11113 361280 140772 361328
rect 426832 361372 434038 361482
rect 11113 336620 11702 361280
rect 15816 358120 16116 361280
rect 426832 360352 427014 361372
rect 433904 361243 434038 361372
rect 433904 361187 581287 361243
rect 433904 360563 580208 361187
rect 581211 360563 581287 361187
rect 433904 360507 581287 360563
rect 433904 360352 434038 360507
rect 426832 360218 434038 360352
rect 575087 358081 576450 358087
rect 452190 358018 576452 358081
rect 452190 358012 575167 358018
rect 452190 357386 452253 358012
rect 456061 357386 575167 358012
rect 452190 357360 575167 357386
rect 576400 357360 576452 358018
rect 452190 357300 576452 357360
rect 575087 357299 576450 357300
rect 444232 356155 576388 356208
rect 444232 355510 444363 356155
rect 448074 356137 576388 356155
rect 448074 355510 575129 356137
rect 444232 355501 575129 355510
rect 576287 355501 576388 356137
rect 444232 355427 576388 355501
rect 440094 355012 440422 355036
rect 440094 354020 440123 355012
rect 440396 354683 440422 355012
rect 440396 354648 580446 354683
rect 440396 354393 579107 354648
rect 580386 354393 580446 354648
rect 440396 354363 580446 354393
rect 440396 354020 440422 354363
rect 440094 353980 440422 354020
rect 65959 350620 169654 352368
rect 61456 350180 169654 350620
rect 11107 336581 11768 336620
rect 11107 335652 11146 336581
rect 11723 335652 11768 336581
rect 11107 335605 11768 335652
rect 7923 334800 10526 335271
rect 6704 334784 10526 334800
rect 6704 334714 8008 334784
rect 1229 330761 6115 332034
rect 1229 299845 2502 330761
rect 14832 314656 15352 348622
rect 65959 347766 169654 350180
rect 65959 345626 116072 347766
rect 118072 345626 169654 347766
rect 65959 343186 169654 345626
rect 16486 314656 17274 319328
rect 25657 318928 26052 319021
rect 25657 318190 25702 318928
rect 26022 318190 26052 318928
rect 25657 315893 26052 318190
rect 567090 316809 568186 316873
rect 25657 315498 144297 315893
rect 2982 314581 114161 314656
rect 2982 311780 3091 314581
rect 3736 314538 114161 314581
rect 3736 311856 106704 314538
rect 113848 311856 114161 314538
rect 3736 311780 114161 311856
rect 2982 311714 114161 311780
rect 3032 311699 3801 311714
rect 5135 310650 132820 310688
rect 5135 310072 50036 310650
rect 50460 310649 132820 310650
rect 50460 310102 128934 310649
rect 132738 310102 132820 310649
rect 50460 310072 132820 310102
rect 5135 310034 132820 310072
rect 5135 301576 5789 310034
rect 6419 309624 140859 309688
rect 6419 309106 136918 309624
rect 140746 309106 140859 309624
rect 6419 309034 140859 309106
rect 6419 302789 7073 309034
rect 10005 308204 10187 308217
rect 10005 308203 52944 308204
rect 10005 307782 10019 308203
rect 10174 307819 52944 308203
rect 10174 307782 10187 307819
rect 10005 307770 10187 307782
rect 7556 307000 7776 307036
rect 7556 306618 7588 307000
rect 7747 306687 7776 307000
rect 50010 306986 50494 307018
rect 7747 306618 12595 306687
rect 7556 306587 12595 306618
rect 10647 306338 10847 306354
rect 10647 305956 10668 306338
rect 10827 306287 10847 306338
rect 10827 306187 12570 306287
rect 10827 305956 10847 306187
rect 10647 305932 10847 305956
rect 50010 306142 50036 306986
rect 50462 306142 50494 306986
rect 11106 305746 12139 305887
rect 11106 303268 11210 305746
rect 12045 303268 12139 305746
rect 11106 303184 12139 303268
rect 11825 302878 12121 302887
rect 6419 302135 9671 302789
rect 10005 302786 10187 302798
rect 11825 302797 11839 302878
rect 12083 302797 12121 302878
rect 11825 302787 12121 302797
rect 10005 302398 10018 302786
rect 10174 302487 10187 302786
rect 11825 302677 12121 302687
rect 11825 302596 11835 302677
rect 12079 302596 12121 302677
rect 11825 302587 12121 302596
rect 10174 302398 12121 302487
rect 10005 302387 12121 302398
rect 10005 302386 10187 302387
rect 5135 300922 8429 301576
rect 1229 298572 6467 299845
rect 5194 296534 6467 298572
rect 5194 296044 5290 296534
rect 6335 296044 6467 296534
rect 5194 287221 6467 296044
rect 7775 292167 8429 300922
rect 9017 301571 9671 302135
rect 11109 302203 12146 302284
rect 9017 300917 10426 301571
rect 9772 293093 10426 300917
rect 11109 300132 11210 302203
rect 12031 300132 12146 302203
rect 11109 299985 12146 300132
rect 50010 299887 50494 306142
rect 48688 299787 50494 299887
rect 8863 293051 10426 293093
rect 8863 292471 8908 293051
rect 9750 292471 10426 293051
rect 8863 292434 10426 292471
rect 7037 292119 8429 292167
rect 7037 291597 7102 292119
rect 8352 291597 8429 292119
rect 7037 291557 8429 291597
rect 5194 286612 5242 287221
rect 6400 286612 6467 287221
rect 5194 286492 6467 286612
rect 7775 286306 8429 291557
rect 9775 287991 10426 292434
rect 9775 287428 9820 287991
rect 10389 287428 10426 287991
rect 9775 287372 10426 287428
rect 7775 285650 7809 286306
rect 8396 285650 8429 286306
rect 7775 285622 8429 285650
rect 52471 241286 52944 307819
rect 91077 305694 100259 306338
rect 91077 303297 91244 305694
rect 100075 303297 100259 305694
rect 91077 290368 100259 303297
rect 143902 299188 144297 315498
rect 567090 315844 567177 316809
rect 568123 315844 568186 316809
rect 444188 310336 448173 310483
rect 444188 309389 444353 310336
rect 448020 310314 448173 310336
rect 448020 310201 566355 310314
rect 448020 309466 565640 310201
rect 448020 309389 448173 309466
rect 444188 309275 448173 309389
rect 565507 309073 565640 309466
rect 566219 309073 566355 310201
rect 452182 306969 456175 307051
rect 452182 306064 452287 306969
rect 456063 306815 456175 306969
rect 456063 306470 564765 306815
rect 456063 306178 564258 306470
rect 456063 306064 456175 306178
rect 452182 305976 456175 306064
rect 564128 305360 564258 306178
rect 564610 305360 564765 306470
rect 143902 298793 270114 299188
rect 269719 295188 270114 298793
rect 444174 298616 448176 298680
rect 444174 298374 444258 298616
rect 322545 298085 326987 298248
rect 322545 297074 322695 298085
rect 269719 295162 283999 295188
rect 263426 294796 265741 294863
rect 128541 294713 265741 294796
rect 269719 294793 283572 295162
rect 128541 294706 263662 294713
rect 128541 293979 136946 294706
rect 140744 293984 263662 294706
rect 265591 293984 265741 294713
rect 140744 293979 265741 293984
rect 128541 293892 265741 293979
rect 263426 293791 265741 293892
rect 283533 293605 283572 294793
rect 283964 293605 283999 295162
rect 283533 293564 283999 293605
rect 291775 294833 322695 297074
rect 245574 293196 247889 293256
rect 128541 293106 247904 293196
rect 128541 293105 245788 293106
rect 128541 292378 128935 293105
rect 132733 292378 245788 293105
rect 128541 292377 245788 292378
rect 247717 292377 247904 293106
rect 128541 292292 247904 292377
rect 245574 292184 247889 292292
rect 91077 286830 169654 290368
rect 289080 288789 290237 288826
rect 289080 288764 289130 288789
rect 91077 284192 122182 286830
rect 124562 284192 169654 286830
rect 91077 281186 169654 284192
rect 284823 288524 289130 288764
rect 290210 288524 290237 288789
rect 284823 288517 290237 288524
rect 284823 278813 285070 288517
rect 289080 288488 290237 288517
rect 289072 287302 290229 287341
rect 289072 287288 289114 287302
rect 285228 287041 289114 287288
rect 284759 278775 285073 278813
rect 284759 278144 284796 278775
rect 285034 278144 285073 278775
rect 284759 278096 285073 278144
rect 285228 276725 285475 287041
rect 289072 287037 289114 287041
rect 290194 287037 290229 287302
rect 289072 287003 290229 287037
rect 289065 286661 290222 286695
rect 289065 286650 289110 286661
rect 285677 286403 289110 286650
rect 285142 276685 285477 276725
rect 285142 276044 285179 276685
rect 285438 276044 285477 276685
rect 285142 276002 285477 276044
rect 285677 274561 285924 286403
rect 289065 286396 289110 286403
rect 290190 286396 290222 286661
rect 289065 286357 290222 286396
rect 291775 278473 293460 294833
rect 322546 293780 322695 294833
rect 322545 293607 322695 293780
rect 326820 294787 326987 298085
rect 444172 297974 444258 298374
rect 444174 297698 444258 297974
rect 448110 298374 448176 298616
rect 448110 297974 482216 298374
rect 448110 297698 448176 297974
rect 444174 297624 448176 297698
rect 332132 296686 456374 296787
rect 332132 295951 444240 296686
rect 448055 295951 456374 296686
rect 332132 295883 456374 295951
rect 481816 296272 482216 297974
rect 326820 293883 326989 294787
rect 326820 293607 326987 293883
rect 322545 293467 326987 293607
rect 321062 292959 323381 293065
rect 332132 292959 333036 295883
rect 481816 295872 517992 296272
rect 481816 295774 516181 295812
rect 481816 295445 513273 295774
rect 513751 295445 516181 295774
rect 481816 295412 516181 295445
rect 338902 295187 341217 295247
rect 338887 295119 456374 295187
rect 338887 295097 452291 295119
rect 338887 294368 339074 295097
rect 341003 294384 452291 295097
rect 456106 294384 456374 295119
rect 341003 294368 456374 294384
rect 338887 294283 456374 294368
rect 338902 294175 341217 294283
rect 452178 293534 456176 293586
rect 452178 293258 452238 293534
rect 321062 292916 333036 292959
rect 321062 292187 321212 292916
rect 323141 292187 333036 292916
rect 452176 292858 452238 293258
rect 452178 292590 452238 292858
rect 456120 293258 456176 293534
rect 481816 293258 482216 295412
rect 456120 292858 482216 293258
rect 492058 294952 516181 295352
rect 456120 292590 456176 292858
rect 321062 292055 333036 292187
rect 421275 292454 422943 292553
rect 452178 292534 456176 292590
rect 421275 292142 421370 292454
rect 321062 291994 323381 292055
rect 322557 291992 323381 291994
rect 350141 292005 421370 292142
rect 422855 292005 422943 292454
rect 350141 291994 422943 292005
rect 350141 291254 350289 291994
rect 421275 291915 422943 291994
rect 423790 291865 425460 291985
rect 423790 291656 423897 291865
rect 299742 291106 350289 291254
rect 350938 291416 423897 291656
rect 425382 291416 425460 291865
rect 350938 291344 425460 291416
rect 350938 291343 425047 291344
rect 299742 286011 299890 291106
rect 350938 290698 351251 291343
rect 300298 290385 351251 290698
rect 300298 286012 300611 290385
rect 492058 290324 492458 294952
rect 493574 294492 516181 294892
rect 417050 287604 492543 290324
rect 299307 285969 299931 286011
rect 299307 285048 299365 285969
rect 299882 285048 299931 285969
rect 299307 284990 299931 285048
rect 300260 285959 300884 286012
rect 300260 285038 300312 285959
rect 300829 285038 300884 285959
rect 300260 284991 300884 285038
rect 307850 284381 313094 284382
rect 293611 284232 313094 284381
rect 293611 282800 306274 284232
rect 312971 282800 313094 284232
rect 293611 282696 313094 282800
rect 417050 284006 427136 287604
rect 430734 284006 492543 287604
rect 293611 278473 295296 282696
rect 417050 281142 492543 284006
rect 466202 279504 473690 279505
rect 493574 279504 493974 294492
rect 495026 283932 495434 283962
rect 495026 283618 495054 283932
rect 495406 283618 495434 283932
rect 495026 283590 495434 283618
rect 466202 279404 493974 279504
rect 466202 278013 466365 279404
rect 473556 279104 493974 279404
rect 473556 278013 473690 279104
rect 466202 277893 473690 278013
rect 442680 277307 443004 277338
rect 442680 277078 442709 277307
rect 442672 276942 442709 277078
rect 442680 276714 442709 276942
rect 442977 277078 443004 277307
rect 495150 277078 495286 283590
rect 497587 279858 498079 279892
rect 497587 279505 497633 279858
rect 498017 279505 498079 279858
rect 497587 279457 498079 279505
rect 442977 276942 495286 277078
rect 442977 276714 443004 276942
rect 442680 276686 443004 276714
rect 285646 274532 285965 274561
rect 285646 273948 285676 274532
rect 285943 273948 285965 274532
rect 440905 274403 441261 274429
rect 440905 274339 440930 274403
rect 440904 274120 440930 274339
rect 285646 273912 285965 273948
rect 440905 273577 440930 274120
rect 441236 274339 441261 274403
rect 497713 274339 497932 279457
rect 441236 274120 497932 274339
rect 441236 273577 441261 274120
rect 440905 273540 441261 273577
rect 564128 267662 564765 305360
rect 564128 267178 564172 267662
rect 564723 267178 564765 267662
rect 564128 267113 564765 267178
rect 565507 266037 566355 309073
rect 567090 272468 568186 315844
rect 569251 315568 570067 315681
rect 569251 314111 569330 315568
rect 569965 314111 570067 315568
rect 569251 313992 570067 314111
rect 571015 314309 572629 314379
rect 567084 272396 568186 272468
rect 567084 271604 567218 272396
rect 568058 271604 568186 272396
rect 567084 271516 568186 271604
rect 565507 265643 565565 266037
rect 566309 265643 566355 266037
rect 565507 265581 566355 265643
rect 466249 255107 473735 255449
rect 466249 247031 466498 255107
rect 473424 247031 473735 255107
rect 525004 250793 525194 250820
rect 525004 250783 525018 250793
rect 525001 250571 525018 250783
rect 525156 250571 525194 250793
rect 525001 250533 525194 250571
rect 529531 250576 529721 250610
rect 525001 250090 525182 250533
rect 529531 250354 529560 250576
rect 529698 250354 529721 250576
rect 529531 250323 529721 250354
rect 529915 250560 530105 250601
rect 529915 250338 529935 250560
rect 530073 250338 530105 250560
rect 525001 250059 525191 250090
rect 525001 249837 525018 250059
rect 525156 249837 525191 250059
rect 525001 249803 525191 249837
rect 529531 249827 529712 250323
rect 529915 250314 530105 250338
rect 530275 250584 530465 250614
rect 530275 250362 530303 250584
rect 530441 250362 530465 250584
rect 530275 250327 530465 250362
rect 529915 249833 530096 250314
rect 530277 249849 530458 250327
rect 529529 249788 529719 249827
rect 529529 249566 529549 249788
rect 529687 249566 529719 249788
rect 529529 249540 529719 249566
rect 529911 249795 530101 249833
rect 529911 249573 529940 249795
rect 530078 249573 530101 249795
rect 529911 249546 530101 249573
rect 530275 249808 530465 249849
rect 530275 249586 530288 249808
rect 530426 249586 530465 249808
rect 530275 249562 530465 249586
rect 466249 242640 473735 247031
rect 567090 242640 568186 271516
rect 466249 241544 568186 242640
rect 52471 240813 163138 241286
rect 106501 232157 114025 232502
rect 106501 224846 106878 232157
rect 113676 224846 114025 232157
rect 4152 220396 9590 220510
rect 4152 215890 4310 220396
rect 9440 215890 9590 220396
rect 10300 220037 12561 220083
rect 10300 218145 10348 220037
rect 11403 218145 12561 220037
rect 10300 218090 12561 218145
rect 4152 215436 9590 215890
rect 4152 210800 4232 215436
rect 9414 210800 9590 215436
rect 4152 210358 9590 210800
rect 4152 205852 4284 210358
rect 9414 205852 9590 210358
rect 4152 205690 9590 205852
rect 106501 201306 114025 224846
rect 162665 206388 163138 240813
rect 466249 221314 473735 241544
rect 424030 213716 462592 214220
rect 162665 206339 165944 206388
rect 162665 205964 164278 206339
rect 165881 205964 165944 206339
rect 424030 206187 424534 213716
rect 433802 211499 434337 211589
rect 433802 209657 433885 211499
rect 434271 209657 434337 211499
rect 433802 206427 434337 209657
rect 436812 211474 437347 211581
rect 436812 209632 436894 211474
rect 437280 209632 437347 211474
rect 436812 206501 437347 209632
rect 462088 209011 462592 213716
rect 466249 211313 466529 221314
rect 473424 211313 473735 221314
rect 466249 210816 473735 211313
rect 569421 209011 569925 313992
rect 571015 313895 571103 314309
rect 572537 313895 572629 314309
rect 571015 313812 572629 313895
rect 571068 273900 571499 313812
rect 581398 298423 581537 298437
rect 581398 297785 581414 298423
rect 581521 297904 581537 298423
rect 582324 298422 582463 298444
rect 582324 297904 582339 298422
rect 581521 297785 582339 297904
rect 581398 297784 582339 297785
rect 582446 297784 582463 298422
rect 581398 297772 582463 297784
rect 581398 297769 582450 297772
rect 581398 297765 581537 297769
rect 570360 273469 571499 273900
rect 570360 237109 570791 273469
rect 578267 270783 579168 270845
rect 578267 270782 578316 270783
rect 570360 235260 570396 237109
rect 570764 235260 570791 237109
rect 570360 235216 570791 235260
rect 571178 270551 578316 270782
rect 462088 208507 569925 209011
rect 162665 205915 165944 205964
rect 423012 205978 425159 206187
rect 423012 205481 423193 205978
rect 424985 205481 425159 205978
rect 423012 205360 425159 205481
rect 263426 204796 265741 204863
rect 127498 204723 265741 204796
rect 127498 203968 136923 204723
rect 140755 204713 265741 204723
rect 140755 203984 263662 204713
rect 265591 203984 265741 204713
rect 140755 203968 265741 203984
rect 127498 203892 265741 203968
rect 263426 203791 265741 203892
rect 321050 204787 323365 204854
rect 433802 204838 433860 206427
rect 321050 204704 422460 204787
rect 321050 203975 321200 204704
rect 323129 203975 422460 204704
rect 433807 204374 433860 204838
rect 434276 205863 434337 206427
rect 436810 206411 437347 206501
rect 434276 204374 434338 205863
rect 433807 204288 434338 204374
rect 436810 204358 436868 206411
rect 437284 204358 437347 206411
rect 436810 204293 437347 204358
rect 436810 204292 437341 204293
rect 321050 203883 422460 203975
rect 321050 203782 323365 203883
rect 245574 203196 247889 203256
rect 127498 203118 247904 203196
rect 127498 202363 128929 203118
rect 132761 203106 247904 203118
rect 132761 202377 245788 203106
rect 247717 202377 247904 203106
rect 132761 202363 247904 202377
rect 127498 202292 247904 202363
rect 338902 203187 341217 203247
rect 338902 203097 420560 203187
rect 338902 202368 339074 203097
rect 341003 202368 420560 203097
rect 245574 202184 247889 202292
rect 338902 202283 420560 202368
rect 338902 202175 341217 202283
rect 106501 194909 106922 201306
rect 113632 194909 114025 201306
rect 419656 200420 420560 202283
rect 421556 202526 422460 203883
rect 421556 202455 456453 202526
rect 421556 201720 444285 202455
rect 448100 201720 456453 202455
rect 421556 201622 456453 201720
rect 419656 200344 456270 200420
rect 419656 199609 452266 200344
rect 456081 199609 456270 200344
rect 419656 199516 456270 199609
rect 423369 196209 424989 196278
rect 423369 195753 423476 196209
rect 424871 196075 424989 196209
rect 571178 196075 571409 270551
rect 578267 270535 578316 270551
rect 579119 270535 579168 270783
rect 578267 270495 579168 270535
rect 578265 269758 579153 269826
rect 578265 269753 578330 269758
rect 575941 269503 578330 269753
rect 575941 240866 576191 269503
rect 578265 269456 578330 269503
rect 579103 269456 579153 269758
rect 578265 269412 579153 269456
rect 574774 240690 580212 240866
rect 574774 236252 574934 240690
rect 580058 236252 580212 240690
rect 574774 235522 580212 236252
rect 574774 231084 574962 235522
rect 580086 231084 580212 235522
rect 574774 230660 580212 231084
rect 574774 226222 574962 230660
rect 580086 226222 580212 230660
rect 574774 226046 580212 226222
rect 424871 195844 571409 196075
rect 574748 196850 580186 197028
rect 424871 195753 424989 195844
rect 423369 195667 424989 195753
rect 106501 194569 114025 194909
rect 574748 192412 574896 196850
rect 580020 192412 580186 196850
rect 574748 192076 580186 192412
rect 451946 191899 580186 192076
rect 451946 187251 452333 191899
rect 455990 187251 580186 191899
rect 451946 187076 580186 187251
rect 574748 186806 580186 187076
rect 574748 182368 574908 186806
rect 580032 182368 580186 186806
rect 574748 182208 580186 182368
rect 444183 180774 448179 180858
rect 444183 179958 444303 180774
rect 448071 180530 448179 180774
rect 448071 180130 482138 180530
rect 448071 179958 448179 180130
rect 444183 179854 448179 179958
rect 481738 179315 482138 180130
rect 481738 178915 523452 179315
rect 481738 178455 521694 178855
rect 3532 178310 8768 178430
rect 3532 173829 3756 178310
rect 8602 173829 8768 178310
rect 452176 177478 456170 177590
rect 452176 176624 452276 177478
rect 456058 177281 456170 177478
rect 481738 177281 482138 178455
rect 456058 176881 482138 177281
rect 485576 177995 521684 178395
rect 456058 176624 456170 176881
rect 452176 176524 456170 176624
rect 3532 173694 8768 173829
rect 466206 175148 473676 175258
rect 3532 173511 133180 173694
rect 3532 168834 129023 173511
rect 132621 168834 133180 173511
rect 466206 173412 466300 175148
rect 473518 174450 473676 175148
rect 485576 174450 485976 177995
rect 473518 174050 485976 174450
rect 489372 177535 521684 177935
rect 473518 173412 473676 174050
rect 466206 173320 473676 173412
rect 489372 170324 489772 177535
rect 3532 168694 133180 168834
rect 3532 168320 8768 168694
rect 3532 163839 3676 168320
rect 8522 163839 8768 168320
rect 3532 163716 8768 163839
rect 417050 167041 489944 170324
rect 417050 163637 431353 167041
rect 434495 163637 489944 167041
rect 417050 161142 489944 163637
rect 442681 156796 443002 156820
rect 442681 156356 442705 156796
rect 442679 156171 442705 156356
rect 442983 156356 443002 156796
rect 442983 156342 493210 156356
rect 442983 156171 492662 156342
rect 442679 156162 492662 156171
rect 493194 156162 493210 156342
rect 440921 156125 441168 156151
rect 442679 156148 493210 156162
rect 442681 156146 443002 156148
rect 440921 155284 440954 156125
rect 441137 155747 441168 156125
rect 493979 155747 494657 155756
rect 441137 155736 494657 155747
rect 441137 155593 494004 155736
rect 441137 155284 441168 155593
rect 493979 155582 494004 155593
rect 494639 155582 494657 155736
rect 493979 155562 494657 155582
rect 440921 155253 441168 155284
rect 574794 152256 580634 152400
rect 8354 150326 169654 150368
rect 8077 146268 169654 150326
rect 8077 143960 146008 146268
rect 148318 143960 169654 146268
rect 8077 141186 169654 143960
rect 574794 147818 575156 152256
rect 580280 147818 580634 152256
rect 574794 147254 580634 147818
rect 574794 142816 575132 147254
rect 580256 142816 580634 147254
rect 574794 142194 580634 142816
rect 4333 138343 6731 138451
rect 4331 138293 6746 138343
rect 4331 132170 4491 138293
rect 6606 132170 6746 138293
rect 4331 107789 6746 132170
rect 8077 113162 10345 141186
rect 574794 137756 575102 142194
rect 580226 137756 580634 142194
rect 574794 137630 580634 137756
rect 122014 117189 166294 117233
rect 122014 116572 122080 117189
rect 124173 117154 166294 117189
rect 124173 116604 164579 117154
rect 166211 116604 166294 117154
rect 124173 116572 166294 116604
rect 122014 116519 166294 116572
rect 263426 114796 265741 114863
rect 127952 114737 265741 114796
rect 127952 113982 136938 114737
rect 140770 114713 265741 114737
rect 140770 113984 263662 114713
rect 265591 113984 265741 114713
rect 140770 113982 265741 113984
rect 127952 113892 265741 113982
rect 263426 113791 265741 113892
rect 321050 114787 323365 114854
rect 321050 114711 456361 114787
rect 321050 114704 444260 114711
rect 321050 113975 321200 114704
rect 323129 113976 444260 114704
rect 448075 113976 456361 114711
rect 323129 113975 456361 113976
rect 321050 113883 456361 113975
rect 321050 113782 323365 113883
rect 245574 113196 247889 113256
rect 8077 109813 8320 113162
rect 10127 109813 10345 113162
rect 127952 113106 247904 113196
rect 338902 113187 341217 113247
rect 127952 112351 128914 113106
rect 132746 112377 245788 113106
rect 247717 112377 247904 113106
rect 132746 112351 247904 112377
rect 127952 112292 247904 112351
rect 338887 113100 456361 113187
rect 338887 113097 452266 113100
rect 338887 112368 339074 113097
rect 341003 112368 452266 113097
rect 338887 112365 452266 112368
rect 456081 112365 456361 113100
rect 245574 112184 247889 112292
rect 338887 112283 456361 112365
rect 338902 112175 341217 112283
rect 8077 109555 10345 109813
rect 4331 104052 4550 107789
rect 6568 104052 6746 107789
rect 4331 103820 6746 104052
rect 444175 92247 448174 92351
rect 444175 91356 444290 92247
rect 448055 92019 448174 92247
rect 448055 91619 487574 92019
rect 448055 91356 448174 91619
rect 444175 91248 448174 91356
rect 487174 90694 487574 91619
rect 487104 90294 516122 90694
rect 487104 89834 516501 90234
rect 452177 89388 456180 89459
rect 452177 89142 452241 89388
rect 452171 88742 452241 89142
rect 452177 88492 452241 88742
rect 456105 89142 456180 89388
rect 487104 89142 487504 89834
rect 456105 88742 487504 89142
rect 495364 89374 516501 89774
rect 456105 88492 456180 88742
rect 452177 88434 456180 88492
rect 106534 87962 114014 88209
rect 106534 87732 106781 87962
rect 3859 86858 106781 87732
rect 113786 87732 114014 87962
rect 113786 86858 114051 87732
rect 3859 86630 114051 86858
rect 3859 79506 4961 86630
rect 7419 85335 132969 85421
rect 7419 85317 128916 85335
rect 7419 84414 7550 85317
rect 11060 84414 128916 85317
rect 7419 84353 128916 84414
rect 132725 84353 132969 85335
rect 7419 84273 132969 84353
rect 5652 83186 140902 83268
rect 5652 83143 136942 83186
rect 5652 82240 5768 83143
rect 9278 82240 136942 83143
rect 5652 82204 136942 82240
rect 140751 82204 140902 83186
rect 5652 82120 140902 82204
rect 150790 80603 158018 80784
rect 150790 80295 151028 80603
rect 3859 78534 3917 79506
rect 4887 78534 4961 79506
rect 3859 78471 4961 78534
rect 5797 78823 151028 80295
rect 5797 45170 7269 78823
rect 150790 78588 151028 78823
rect 157755 78588 158018 80603
rect 150790 78317 158018 78588
rect 442643 78912 443060 78961
rect 442643 77894 442690 78912
rect 443023 78236 443060 78912
rect 443023 78206 489758 78236
rect 443023 77954 488864 78206
rect 489714 77954 489758 78206
rect 443023 77922 489758 77954
rect 443023 77894 443060 77922
rect 442643 77852 443060 77894
rect 440169 74403 440421 74427
rect 440169 73811 440192 74403
rect 440394 74192 440421 74403
rect 488770 74217 489966 74243
rect 488770 74192 488810 74217
rect 440394 73992 488810 74192
rect 440394 73811 440421 73992
rect 488770 73965 488810 73992
rect 489925 73965 489966 74217
rect 488770 73936 489966 73965
rect 440169 73781 440421 73811
rect 148532 70280 169654 70368
rect 495364 70324 495764 89374
rect 498066 88914 516501 89314
rect 146751 66158 169654 70280
rect 146751 63802 159964 66158
rect 162104 63802 169654 66158
rect 146751 61186 169654 63802
rect 417050 67289 496013 70324
rect 417050 63691 436136 67289
rect 439734 63691 496013 67289
rect 80484 56959 132866 57085
rect 80484 53284 128967 56959
rect 132708 53284 132866 56959
rect 80484 53164 132866 53284
rect 146751 46454 149672 61186
rect 417050 61142 496013 63691
rect 466219 59292 473683 59375
rect 466219 58179 466321 59292
rect 473542 58976 473683 59292
rect 498066 58976 498466 88914
rect 473542 58576 498466 58976
rect 473542 58179 473683 58576
rect 466219 58099 473683 58179
rect 5820 39493 6396 45170
rect 81943 43276 149672 46454
rect 56490 42522 57962 42524
rect 78726 42317 149672 43276
rect 136362 40865 167859 41116
rect 5652 39422 6511 39493
rect 5652 38923 5712 39422
rect 6434 38923 6511 39422
rect 5652 38883 6511 38923
rect 136362 32718 137083 40865
rect 113034 32468 137083 32718
rect 113034 31500 113278 32468
rect 118898 31547 137083 32468
rect 140503 31610 157632 40865
rect 167451 31610 167859 40865
rect 426799 39173 434047 39338
rect 140503 31547 167859 31610
rect 118898 31500 167859 31547
rect 113034 31270 167859 31500
rect 136362 31139 167859 31270
rect 128832 28804 280822 28976
rect 128832 23480 129020 28804
rect 132614 28758 280822 28804
rect 132614 23492 273418 28758
rect 280424 23492 280822 28758
rect 132614 23480 280822 23492
rect 128832 23252 280822 23480
rect 291775 24480 293460 32589
rect 293611 27790 295296 32589
rect 426799 32240 426979 39173
rect 433851 32240 434047 39173
rect 426799 32090 434047 32240
rect 293611 27651 313157 27790
rect 293611 26209 306753 27651
rect 313014 26209 313157 27651
rect 293611 26105 313157 26209
rect 428910 24480 430595 32090
rect 291775 22795 430595 24480
rect 3527 18165 291000 18190
rect 3527 18157 290103 18165
rect 3527 17264 3562 18157
rect 4344 17264 290103 18157
rect 3527 17259 290103 17264
rect 290967 17259 291000 18165
rect 3527 17232 291000 17259
<< via4 >>
rect 516456 693856 520966 698932
rect 466468 569837 473449 577278
rect 4066 555362 9170 560048
rect 466599 553646 473439 560021
rect 466547 523885 473413 530621
rect 575622 546532 580746 550970
rect 572241 527565 574152 529912
rect 106611 470309 113894 475380
rect 273494 472164 280502 475224
rect 150899 461395 157916 462824
rect 106619 454319 113903 455661
rect 106630 440408 113902 441575
rect 150941 439040 157881 440395
rect 466355 410038 473541 412620
rect 163821 391614 167356 400684
rect 106648 387014 113913 387634
rect 150869 380153 157943 381083
rect 150962 366820 157821 369602
rect 466376 367103 473507 368377
rect 427014 360352 433904 361372
rect 106704 311856 113848 314538
rect 11210 303268 12045 305746
rect 11210 300132 12031 302203
rect 91244 303297 100075 305694
rect 322695 293607 326820 298085
rect 306274 282800 312971 284232
rect 466365 278013 473556 279404
rect 466498 247031 473424 255107
rect 106878 224846 113676 232157
rect 4232 210800 9414 215436
rect 466529 211313 473424 221314
rect 570396 235260 570764 237109
rect 106922 194909 113632 201306
rect 574962 231084 580086 235522
rect 466300 173412 473518 175148
rect 575132 142816 580256 147254
rect 4491 132170 6606 138293
rect 106781 86858 113786 87962
rect 151028 78588 157755 80603
rect 466321 58179 473542 59292
rect 157632 31610 167451 40865
rect 273418 23492 280424 28758
rect 426979 32240 433851 39173
rect 306753 26209 313014 27651
<< metal5 >>
rect 166394 703100 171394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 330094 703100 335094 704800
rect 516238 698932 521238 699090
rect 516238 696670 516456 698932
rect 515321 693856 516456 696670
rect 520966 696670 521238 698932
rect 520966 693856 522787 696670
rect 515321 672866 522787 693856
rect 106520 665257 280703 672722
rect 106520 561595 114019 665257
rect 6412 560186 114019 561595
rect 3942 560048 114019 560186
rect 3942 555362 4066 560048
rect 9170 555362 114019 560048
rect 3942 555186 114019 555362
rect 6412 554130 114019 555186
rect 106520 475380 114019 554130
rect 106520 470309 106611 475380
rect 113894 470309 114019 475380
rect 106520 455661 114019 470309
rect 106520 454319 106619 455661
rect 113903 454319 114019 455661
rect 106520 441575 114019 454319
rect 106520 440408 106630 441575
rect 113902 440408 114019 441575
rect 106520 387634 114019 440408
rect 106520 387014 106648 387634
rect 113913 387014 114019 387634
rect 106520 314538 114019 387014
rect 106520 311856 106704 314538
rect 113848 311856 114019 314538
rect 11007 305746 100229 305828
rect 11007 303268 11210 305746
rect 12045 305694 100229 305746
rect 12045 303297 91244 305694
rect 100075 303297 100229 305694
rect 12045 303268 100229 303297
rect 11007 303187 100229 303268
rect 106520 302347 114019 311856
rect 11007 302203 114019 302347
rect 11007 300132 11210 302203
rect 12031 300132 114019 302203
rect 11007 299886 114019 300132
rect 106520 232157 114019 299886
rect 106520 224846 106878 232157
rect 113676 224846 114019 232157
rect 106520 224434 114019 224846
rect 150783 572691 172377 579941
rect 150783 489095 158033 572691
rect 150783 481845 169318 489095
rect 273238 488701 280703 665257
rect 305969 665400 522787 672866
rect 150783 462824 158033 481845
rect 273238 481236 293998 488701
rect 150783 461395 150899 462824
rect 157916 461395 158033 462824
rect 150783 440395 158033 461395
rect 150783 439040 150941 440395
rect 157881 439040 158033 440395
rect 150783 381083 158033 439040
rect 273238 475224 280703 475600
rect 273238 472164 273494 475224
rect 280502 472164 280703 475224
rect 163332 400684 168774 401219
rect 163332 391614 163821 400684
rect 167356 391614 168774 400684
rect 163332 391172 168774 391614
rect 273238 391276 280703 472164
rect 286533 381833 293998 481236
rect 150783 380153 150869 381083
rect 157943 380153 158033 381083
rect 273240 380558 293998 381833
rect 150783 369602 158033 380153
rect 150783 366820 150962 369602
rect 157821 366820 158033 369602
rect 150783 309095 158033 366820
rect 273238 374368 293998 380558
rect 150783 301845 169318 309095
rect 150783 219095 158033 301845
rect 150783 216733 169318 219095
rect 8595 215634 169318 216733
rect 4098 215436 169318 215634
rect 4098 210800 4232 215436
rect 9414 211845 169318 215436
rect 9414 210800 158033 211845
rect 4098 210634 158033 210800
rect 8595 209483 158033 210634
rect 106520 201306 114019 201663
rect 106520 194909 106922 201306
rect 113632 194909 114019 201306
rect 106520 138452 114019 194909
rect 4506 138451 114019 138452
rect 4333 138293 114019 138451
rect 4333 132170 4491 138293
rect 6606 132170 114019 138293
rect 4333 131986 114019 132170
rect 4333 131971 6731 131986
rect 106520 87962 114019 131986
rect 106520 86858 106781 87962
rect 113786 86858 114019 87962
rect 106520 85771 114019 86858
rect 150783 129095 158033 209483
rect 150783 121845 169318 129095
rect 150783 80603 158033 121845
rect 273238 120698 280703 374368
rect 305969 284232 313435 665400
rect 418431 572089 434054 579339
rect 426804 546276 434054 572089
rect 466215 577278 473681 665400
rect 466215 569837 466468 577278
rect 473449 569837 473681 577278
rect 466215 560021 473681 569837
rect 466215 553646 466599 560021
rect 473439 553646 473681 560021
rect 466215 553211 473681 553646
rect 553960 551280 577018 551988
rect 553960 550970 580932 551280
rect 553960 546532 575622 550970
rect 580746 546532 580932 550970
rect 553960 546280 580932 546532
rect 553960 546276 577018 546280
rect 426804 544738 577018 546276
rect 426804 539026 561210 544738
rect 426804 489339 434054 539026
rect 418431 482089 434054 489339
rect 426804 430706 434054 482089
rect 426216 427736 434054 430706
rect 426804 399339 434054 427736
rect 466215 530621 473681 530943
rect 466215 523885 466547 530621
rect 473413 530016 473681 530621
rect 473413 529912 574258 530016
rect 473413 527565 572241 529912
rect 574152 527565 574258 529912
rect 473413 527489 574258 527565
rect 473413 523885 473681 527489
rect 466215 412769 473681 523885
rect 466206 412620 473703 412769
rect 466206 410038 466355 412620
rect 473541 410038 473703 412620
rect 466206 409865 473703 410038
rect 418431 392089 434054 399339
rect 426804 361372 434054 392089
rect 426804 360352 427014 361372
rect 433904 360352 434054 361372
rect 426804 309339 434054 360352
rect 418431 302089 434054 309339
rect 426804 298253 434054 302089
rect 322531 298085 434054 298253
rect 322531 293607 322695 298085
rect 326820 293607 434054 298085
rect 322531 293461 434054 293607
rect 305969 282800 306274 284232
rect 312971 282800 313435 284232
rect 150783 78588 151028 80603
rect 157755 78588 158033 80603
rect 150783 77477 158033 78588
rect 157255 40865 168455 41208
rect 157255 31610 157632 40865
rect 167451 31610 168455 40865
rect 157255 31208 168455 31610
rect 273238 28758 280703 111386
rect 273238 23492 273418 28758
rect 280424 23492 280703 28758
rect 273238 23034 280703 23492
rect 305969 27651 313435 282800
rect 426804 237151 434054 293461
rect 466215 368506 473681 409865
rect 466215 368377 473688 368506
rect 466215 367103 466376 368377
rect 473507 367103 473688 368377
rect 466215 366922 473688 367103
rect 466215 279404 473681 366922
rect 466215 278013 466365 279404
rect 473556 278013 473681 279404
rect 466215 255107 473681 278013
rect 466215 247031 466498 255107
rect 473424 247031 473681 255107
rect 466215 246663 473681 247031
rect 426804 237109 577018 237151
rect 426804 235260 570396 237109
rect 570764 235850 577018 237109
rect 570764 235522 580166 235850
rect 570764 235260 574962 235522
rect 426804 231084 574962 235260
rect 580086 231084 580166 235522
rect 426804 230850 580166 231084
rect 426804 229901 577018 230850
rect 426804 219339 434054 229901
rect 418431 212089 434054 219339
rect 426804 129339 434054 212089
rect 418431 122089 434054 129339
rect 426804 39339 434054 122089
rect 418431 39173 434054 39339
rect 418431 32240 426979 39173
rect 433851 32240 434054 39173
rect 418431 32089 434054 32240
rect 466215 221314 473681 221672
rect 466215 211313 466529 221314
rect 473424 211313 473681 221314
rect 466215 175148 473681 211313
rect 466215 173412 466300 175148
rect 473518 173412 473681 175148
rect 466215 103777 473681 173412
rect 573526 149883 580992 153349
rect 573534 147254 580992 149883
rect 573534 142816 575132 147254
rect 580256 142816 580992 147254
rect 573534 139533 580992 142816
rect 573526 103777 580992 139533
rect 466215 96311 580992 103777
rect 466215 59292 473681 96311
rect 466215 58179 466321 59292
rect 473542 58179 473681 59292
rect 305969 26209 306753 27651
rect 313014 26209 313435 27651
rect 305969 26129 313435 26209
rect 466215 26129 473681 58179
rect 305969 18663 473687 26129
<< fillblock >>
rect 287497 306699 302657 310031
rect 290225 302778 296473 306103
<< comment >>
rect 0 704800 585600 705600
rect 0 800 800 704800
rect 32567 595771 73552 604698
rect 533438 596264 551793 600607
rect 27798 503403 49688 511786
rect 490101 475858 531086 484785
rect 18736 437627 38275 444818
rect 533336 425671 556320 432270
rect 555953 362177 575334 365076
rect 65678 334437 80405 337219
rect 490913 331801 531898 340728
rect 505488 270377 512694 273447
rect 55520 259233 77588 264983
rect 528454 124046 542202 127516
rect 31573 116309 49227 121391
rect 41661 60172 59315 65254
rect 494643 49119 509259 52791
rect 584800 800 585600 704800
rect 0 0 585600 800
use analog_mux_sel1v8  analog_mux_sel1v8_0
timestamp 1714180253
transform 0 -1 583347 1 0 361407
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_1
timestamp 1714180253
transform 0 1 5348 1 0 462156
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_2
timestamp 1714180253
transform -1 0 6199 0 1 427752
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_3
timestamp 1714180253
transform 0 1 3252 1 0 296809
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_4
timestamp 1714180253
transform 0 1 2828 1 0 339990
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_5
timestamp 1714180253
transform 0 1 3477 1 0 39710
box -5530 -288 4452 6736
use bias_generator  bias_generator_0
timestamp 1714594028
transform 0 -1 291742 1 0 33373
box -1132 -6353 249191 3114
use font_4C  font_4C_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766404
transform 1 0 295208 0 1 307055
box 0 0 1080 2520
use font_4F  font_4F_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598767855
transform 1 0 296660 0 1 307074
box 0 0 1080 2520
use font_4F  font_4F_1
timestamp 1598767855
transform 1 0 298113 0 1 307092
box 0 0 1080 2520
use font_5A  font_5A_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598772956
transform 1 0 299565 0 1 307111
box 0 0 1080 2520
use font_30  font_30_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786981
transform 1 0 292120 0 1 303139
box 0 0 1080 2520
use font_32  font_32_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787041
transform 1 0 290686 0 1 303118
box 0 0 1080 2520
use font_32  font_32_1
timestamp 1598787041
transform 1 0 293535 0 1 303118
box 0 0 1080 2520
use font_34  font_34_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787136
transform 1 0 295024 0 1 303154
box 0 0 1080 2520
use font_41  font_41_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763107
transform 1 0 293756 0 1 307074
box 0 0 1080 2520
use font_41  font_41_1
timestamp 1598763107
transform 1 0 300982 0 1 307129
box 0 0 1080 2520
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 287836 0 1 307088
box 0 0 1080 2520
use font_48  font_48_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765560
transform 1 0 289326 0 1 307111
box 0 0 1080 2520
use font_49  font_49_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765816
transform 1 0 290833 0 1 307111
box 0 0 1080 2520
use font_50  font_50_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768087
transform 1 0 292285 0 1 307092
box 0 0 1080 2520
use isolated_switch_ena1v8  isolated_switch_ena1v8_0
timestamp 1714180201
transform 1 0 579104 0 -1 497212
box 0 0 4162 6736
use isolated_switch_ena1v8  isolated_switch_ena1v8_1
timestamp 1714180201
transform 1 0 579484 0 -1 272314
box 0 0 4162 6736
use isolated_switch_ena1v8  isolated_switch_ena1v8_2
timestamp 1714180201
transform 1 0 573106 0 -1 316768
box 0 0 4162 6736
use isolated_switch_ena1v8  isolated_switch_ena1v8_4
timestamp 1714180201
transform 1 0 579514 0 -1 586638
box 0 0 4162 6736
use isolated_switch_ena1v8  isolated_switch_ena1v8_5
timestamp 1714180201
transform -1 0 7186 0 -1 384878
box 0 0 4162 6736
use sky130_rodovalho_ip__lpopamp  lpopamp_0 ../dependencies//sky130_rodovalho_ip__lpopamp/mag
timestamp 1714587215
transform 0 -1 48697 -1 0 299887
box -7000 0 81800 36580
use lvl_shift_invert  lvl_shift_invert_0
timestamp 1714065493
transform 0 -1 14197 1 0 286759
box -2394 4352 3500 6736
use power_stage  power_stage_0
array 0 6 90000 0 0 -111006
timestamp 1714671808
transform 0 -1 234941 1 0 120408
box -89200 -44204 -9499 66802
use power_stage  power_stage_1
array 0 6 90000 0 0 111006
timestamp 1714671808
transform 0 1 351850 1 0 120408
box -89200 -44204 -9499 66802
use sky130_ajc_ip__brownout  sky130_ajc_ip__brownout_0 ../dependencies//sky130_ajc_ip__brownout/mag
timestamp 1713419710
transform 0 -1 557384 -1 0 89090
box -1604 -1987 43293 41283
use sky130_ajc_ip__overvoltage  sky130_ajc_ip__overvoltage_0 ../dependencies//sky130_ajc_ip__overvoltage/mag
timestamp 1713210720
transform 0 -1 550164 -1 0 176882
box -2433 -2390 42464 28880
use sky130_ajc_ip__por  sky130_ajc_ip__por_0 ../dependencies//sky130_ajc_ip__por/mag
timestamp 1713454396
transform 0 -1 557064 -1 0 294668
box -1604 -1987 43293 41283
use sky130_ak_ip__comparator  sky130_ak_ip__comparator_0 ../dependencies//sky130_ak_ip__comparator/mag
timestamp 1714760001
transform 0 -1 28376 1 0 319360
box -1900 -33700 39700 13700
use sky130_be_ip__lsxo  sky130_be_ip__lsxo_0 ../dependencies//sky130_be_ip__lsxo/mag
timestamp 1714591373
transform 0 -1 558491 1 0 410746
box 1476 -23704 25570 -812
use sky130_cw_ip__bandgap  sky130_cw_ip__bandgap_0 ../dependencies//sky130_cw_ip/mag
timestamp 1715026686
transform 1 0 38648 0 1 42266
box -5734 12 42048 14837
use sky130_ht_ip__hsxo_cpz1  sky130_ht_ip__hsxo_cpz1_0 ../dependencies//sky130_ht_ip__hsxo_cpz1/mag
timestamp 1714659811
transform 1 0 13043 0 1 95673
box -3162 -7320 32492 17749
use sky130_od_ip__tempsensor_ext_vp  sky130_od_ip__tempsensor_ext_vp_0 ../dependencies//sky130_od_ip__tempsensor/mag
timestamp 1713856378
transform 1 0 9095 0 1 442073
box -584 -5030 6610 3202
use sky130_td_ip__opamp_hp  sky130_td_ip__opamp_hp_0 ../dependencies//sky130_td_ip__opamp_hp/mag
timestamp 1714591961
transform 0 1 10847 1 0 489761
box -7724 -6929 51340 16206
use sky130_vbl_ip__overvoltage  sky130_vbl_ip__overvoltage_0 ../dependencies//sky130_vbl_ip__overvoltage/mag
timestamp 1714660490
transform 1 0 539503 0 1 576713
box -18218 -4002 24405 17489
<< labels >>
flabel metal4 15162 171077 15162 171077 0 FreeSans 16000 0 0 0 vssd2
flabel metal4 13496 642110 13496 642110 0 FreeSans 16000 0 0 0 vccd2
flabel comment 542585 598389 542585 598389 0 FreeSans 16000 0 0 0 overvoltage
flabel comment 544548 428758 544548 428758 0 FreeSans 16000 0 0 0 LSXO
flabel metal4 26979 17673 26979 17673 0 FreeSans 16000 0 0 0 bias_reference_voltage
flabel comment 29461 503602 46827 511520 0 FreeSans 16000 0 0 0 HGBW_op_amp
flabel comment 29455 441019 29455 441019 0 FreeSans 16000 0 0 0 temp_sensor
flabel comment 66756 261907 66756 261907 0 FreeSans 16000 0 0 0 LP_op_amp
flabel comment 73088 335906 73088 335906 0 FreeSans 16000 0 0 0 comparator
flabel comment 40401 118985 40401 118985 0 FreeSans 16000 180 0 0 HSXO
flabel comment 535328 125714 535328 125714 0 FreeSans 16000 180 0 0 overvoltage
flabel comment 565437 363854 565447 363854 0 FreeSans 16000 0 0 0 1.2V_reference
flabel comment 509358 271777 509358 271777 0 FreeSans 16000 180 0 0 por
flabel comment 51234 600438 51234 600438 0 FreeSans 16000 0 0 0 this_space_for_rent
flabel comment 508768 480525 508768 480525 0 FreeSans 16000 0 0 0 this_space_for_rent
flabel comment 509580 336468 509580 336468 0 FreeSans 16000 0 0 0 this_space_for_rent
flabel comment 502185 50921 502185 50921 0 FreeSans 16000 180 0 0 brownout
flabel metal2 s 180988 0 181100 1280 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 184534 0 184646 1280 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 195172 0 195284 1280 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 198718 0 198830 1280 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 202264 0 202376 1280 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205810 0 205922 1280 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 209356 0 209468 1280 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 216448 0 216560 1280 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219994 0 220106 1280 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 223540 0 223652 1280 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 227086 0 227198 1280 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 230632 0 230744 1280 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 234178 0 234290 1280 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 237724 0 237836 1280 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 241270 0 241382 1280 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244816 0 244928 1280 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 248362 0 248474 1280 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251908 0 252020 1280 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 255454 0 255566 1280 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 259000 0 259112 1280 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 262546 0 262658 1280 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 266092 0 266204 1280 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 269638 0 269750 1280 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 273184 0 273296 1280 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 276730 0 276842 1280 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 280276 0 280388 1280 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283822 0 283934 1280 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 287368 0 287480 1280 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290914 0 291026 1280 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 294460 0 294572 1280 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 298006 0 298118 1280 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 301552 0 301664 1280 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 305098 0 305210 1280 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 312190 0 312302 1280 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 319282 0 319394 1280 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 326374 0 326486 1280 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329920 0 330032 1280 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 333466 0 333578 1280 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 337012 0 337124 1280 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 340558 0 340670 1280 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 344104 0 344216 1280 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 347650 0 347762 1280 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 358288 0 358400 1280 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361834 0 361946 1280 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 365380 0 365492 1280 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368926 0 369038 1280 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 372472 0 372584 1280 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 376018 0 376130 1280 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 379564 0 379676 1280 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 383110 0 383222 1280 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 386656 0 386768 1280 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 390202 0 390314 1280 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 393748 0 393860 1280 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 397294 0 397406 1280 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400840 0 400952 1280 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 404386 0 404498 1280 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407932 0 408044 1280 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 411478 0 411590 1280 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 415024 0 415136 1280 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 418570 0 418682 1280 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 422116 0 422228 1280 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 425662 0 425774 1280 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 429208 0 429320 1280 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 432754 0 432866 1280 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 436300 0 436412 1280 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439846 0 439958 1280 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 443392 0 443504 1280 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 446938 0 447050 1280 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 450484 0 450596 1280 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 454030 0 454142 1280 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 457576 0 457688 1280 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 461122 0 461234 1280 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 464668 0 464780 1280 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 468214 0 468326 1280 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 471760 0 471872 1280 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 475306 0 475418 1280 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478852 0 478964 1280 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 482398 0 482510 1280 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485944 0 486056 1280 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 489490 0 489602 1280 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 493036 0 493148 1280 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 496582 0 496694 1280 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 500128 0 500240 1280 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 503674 0 503786 1280 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 507220 0 507332 1280 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 510766 0 510878 1280 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 514312 0 514424 1280 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 517858 0 517970 1280 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 521404 0 521516 1280 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524950 0 525062 1280 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 528496 0 528608 1280 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 532042 0 532154 1280 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 535588 0 535700 1280 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 539134 0 539246 1280 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541498 0 541610 1280 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 548590 0 548702 1280 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 552136 0 552248 1280 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 556864 0 556976 1280 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 560410 0 560522 1280 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563956 0 564068 1280 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 567502 0 567614 1280 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal3 s 583100 678784 585600 683784 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 584320 590272 585600 590384 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s 584320 589090 585600 589202 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s 584320 584362 585600 584474 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s 584320 500850 585600 500962 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 584320 499668 585600 499780 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 584320 494940 585600 495052 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 584320 451700 585600 451812 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 584320 407278 585600 407390 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 584320 360856 585600 360968 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 584320 314452 585600 314564 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 584320 275940 585600 276052 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 584320 274758 585600 274870 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 584320 270030 585600 270142 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s 584320 95918 585600 96030 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 584320 94736 585600 94848 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 584320 51260 585600 51372 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 584320 50078 585600 50190 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 584320 24802 585600 24914 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 584320 23620 585600 23732 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 584320 20074 585600 20186 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 584320 18892 585600 19004 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 584320 15346 585600 15458 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 584320 14164 585600 14276 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 584320 10618 585600 10730 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s 584320 9436 585600 9548 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s 584320 5890 585600 6002 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 584320 320362 585600 320474 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 584320 319180 585600 319292 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 584320 4708 585600 4820 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 800 163688 2460 168488 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal3 s 800 550242 2460 555042 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 800 205688 2460 210488 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 800 634642 2460 639442 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 567394 703100 572394 705600 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 521394 703140 526194 705600 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 511394 703140 516194 705600 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 466194 703100 471194 705600 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 414194 703100 419194 705600 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 330094 703100 335094 705600 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 218094 703100 223094 705600 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 166394 703100 171394 705600 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 120994 703100 125994 705600 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68994 703100 73994 705600 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16994 703100 21994 705600 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 800 681042 2500 686042 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 800 644642 2460 649442 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 800 560242 2460 565042 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 511148 1280 511260 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s 0 469108 1280 469220 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s 0 425886 1280 425998 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 0 382664 1280 382776 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 0 377936 1280 378048 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s 0 376754 1280 376866 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s 0 339442 1280 339554 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s 0 296220 1280 296332 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s 0 253198 1280 253310 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s 800 215688 2460 220488 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 800 173688 2460 178488 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 125576 1280 125688 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s 0 82354 1280 82466 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s 0 39132 1280 39244 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s 0 34404 1280 34516 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s 0 33222 1280 33334 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s 0 17710 1280 17822 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 0 12982 1280 13094 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s 0 11800 1280 11912 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s 0 8254 1280 8366 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s 0 7072 1280 7184 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s 583140 137630 585600 142430 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 583140 182230 585600 187030 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 583140 226030 585600 230830 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 583140 541362 585600 546162 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 583140 630584 585600 635384 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal2 s 571048 0 571160 1280 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 191626 0 191738 1280 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 188080 0 188192 1280 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 131344 0 131456 1280 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 134890 0 135002 1280 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 138436 0 138548 1280 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 141982 0 142094 1280 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 145528 0 145640 1280 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 149074 0 149186 1280 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 152620 0 152732 1280 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 156166 0 156278 1280 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 159712 0 159824 1280 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 163258 0 163370 1280 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 166804 0 166916 1280 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 170350 0 170462 1280 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173896 0 174008 1280 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 177442 0 177554 1280 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel comment 50489 62848 50489 62848 0 FreeSans 16000 180 0 0 bandgap
flabel metal2 s 546226 0 546338 1280 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal3 s 0 2344 1280 2456 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 0 3526 1280 3638 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 0 16528 1280 16640 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 0 37950 1280 38062 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s 0 81172 1280 81284 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s 0 76444 1280 76556 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s 0 77626 1280 77738 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s 0 119666 1280 119778 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s 0 120848 1280 120960 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s 0 124394 1280 124506 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s 0 247288 1280 247400 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s 0 248470 1280 248582 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s 0 252016 1280 252128 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s 0 290310 1280 290422 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 0 291492 1280 291604 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 0 295038 1280 295150 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s 0 333532 1280 333644 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s 0 334714 1280 334826 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s 0 338260 1280 338372 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s 0 381482 1280 381594 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s 0 419976 1280 420088 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s 0 421158 1280 421270 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s 0 424704 1280 424816 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 0 463198 1280 463310 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s 0 464380 1280 464492 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s 0 467926 1280 468038 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s 0 506420 1280 506532 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s 0 507602 1280 507714 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s 0 512330 1280 512442 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s 584320 271212 585600 271324 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s 584320 315634 585600 315746 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 584320 359674 585600 359786 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 584320 364402 585600 364514 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal3 s 584320 365584 585600 365696 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 584320 406096 585600 406208 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 584320 410824 585600 410936 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 584320 412006 585600 412118 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 584320 450518 585600 450630 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 584320 455246 585600 455358 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 584320 456428 585600 456540 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 584320 496122 585600 496234 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 584320 585544 585600 585656 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal2 s 126616 0 126728 1280 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 127798 0 127910 1280 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 130162 0 130274 1280 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 133708 0 133820 1280 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 137254 0 137366 1280 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 140800 0 140912 1280 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 144346 0 144458 1280 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 147892 0 148004 1280 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 151438 0 151550 1280 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 154984 0 155096 1280 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 158530 0 158642 1280 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 162076 0 162188 1280 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 165622 0 165734 1280 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 169168 0 169280 1280 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 172714 0 172826 1280 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 176260 0 176372 1280 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179806 0 179918 1280 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 183352 0 183464 1280 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186898 0 187010 1280 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 190444 0 190556 1280 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193990 0 194102 1280 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 197536 0 197648 1280 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 201082 0 201194 1280 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 204628 0 204740 1280 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 208174 0 208286 1280 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 211720 0 211832 1280 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 212902 0 213014 1280 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215266 0 215378 1280 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218812 0 218924 1280 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 222358 0 222470 1280 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225904 0 226016 1280 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 229450 0 229562 1280 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 232996 0 233108 1280 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 236542 0 236654 1280 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 240088 0 240200 1280 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 243634 0 243746 1280 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 247180 0 247292 1280 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 250726 0 250838 1280 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 254272 0 254384 1280 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257818 0 257930 1280 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 261364 0 261476 1280 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264910 0 265022 1280 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 268456 0 268568 1280 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 272002 0 272114 1280 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 275548 0 275660 1280 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 279094 0 279206 1280 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 282640 0 282752 1280 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 286186 0 286298 1280 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 289732 0 289844 1280 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 293278 0 293390 1280 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296824 0 296936 1280 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 300370 0 300482 1280 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 303916 0 304028 1280 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 307462 0 307574 1280 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 308644 0 308756 1280 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311008 0 311120 1280 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 314554 0 314666 1280 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 315736 0 315848 1280 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318100 0 318212 1280 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 321646 0 321758 1280 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 322828 0 322940 1280 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325192 0 325304 1280 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 328738 0 328850 1280 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 332284 0 332396 1280 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335830 0 335942 1280 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 339376 0 339488 1280 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342922 0 343034 1280 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 346468 0 346580 1280 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 350014 0 350126 1280 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 353560 0 353672 1280 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 351196 0 351308 1280 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 354742 0 354854 1280 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357106 0 357218 1280 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 360652 0 360764 1280 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 364198 0 364310 1280 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 367744 0 367856 1280 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 371290 0 371402 1280 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 374836 0 374948 1280 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 378382 0 378494 1280 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381928 0 382040 1280 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 385474 0 385586 1280 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 389020 0 389132 1280 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 392566 0 392678 1280 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 396112 0 396224 1280 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 399658 0 399770 1280 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 403204 0 403316 1280 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 406750 0 406862 1280 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 410296 0 410408 1280 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413842 0 413954 1280 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 417388 0 417500 1280 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420934 0 421046 1280 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 424480 0 424592 1280 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 428026 0 428138 1280 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 431572 0 431684 1280 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 435118 0 435230 1280 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 438664 0 438776 1280 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 442210 0 442322 1280 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 445756 0 445868 1280 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 449302 0 449414 1280 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452848 0 452960 1280 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 456394 0 456506 1280 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459940 0 460052 1280 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 463486 0 463598 1280 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 467032 0 467144 1280 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 470578 0 470690 1280 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 474124 0 474236 1280 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 477670 0 477782 1280 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 481216 0 481328 1280 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 484762 0 484874 1280 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 488308 0 488420 1280 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491854 0 491966 1280 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 495400 0 495512 1280 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498946 0 499058 1280 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 502492 0 502604 1280 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 506038 0 506150 1280 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 509584 0 509696 1280 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 513130 0 513242 1280 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 516676 0 516788 1280 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 520222 0 520334 1280 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 523768 0 523880 1280 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 527314 0 527426 1280 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530860 0 530972 1280 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 534406 0 534518 1280 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537952 0 538064 1280 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 542680 0 542792 1280 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545044 0 545156 1280 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 549772 0 549884 1280 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 553318 0 553430 1280 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 555682 0 555794 1280 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 559228 0 559340 1280 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 562774 0 562886 1280 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 566320 0 566432 1280 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569866 0 569978 1280 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 573412 0 573524 1280 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576958 0 577070 1280 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 574594 0 574706 1280 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 578140 0 578252 1280 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
<< end >>
