magic
tech sky130A
magscale 1 2
timestamp 1713888873
<< pwell >>
rect -6758 -3582 6758 3582
<< psubdiff >>
rect -6722 3512 -6626 3546
rect 6626 3512 6722 3546
rect -6722 3450 -6688 3512
rect 6688 3450 6722 3512
rect -6722 -3512 -6688 -3450
rect 6688 -3512 6722 -3450
rect -6722 -3546 -6626 -3512
rect 6626 -3546 6722 -3512
<< psubdiffcont >>
rect -6626 3512 6626 3546
rect -6722 -3450 -6688 3450
rect 6688 -3450 6722 3450
rect -6626 -3546 6626 -3512
<< xpolycontact >>
rect -6592 2984 -6522 3416
rect -6592 -3416 -6522 -2984
rect -6426 2984 -6356 3416
rect -6426 -3416 -6356 -2984
rect -6260 2984 -6190 3416
rect -6260 -3416 -6190 -2984
rect -6094 2984 -6024 3416
rect -6094 -3416 -6024 -2984
rect -5928 2984 -5858 3416
rect -5928 -3416 -5858 -2984
rect -5762 2984 -5692 3416
rect -5762 -3416 -5692 -2984
rect -5596 2984 -5526 3416
rect -5596 -3416 -5526 -2984
rect -5430 2984 -5360 3416
rect -5430 -3416 -5360 -2984
rect -5264 2984 -5194 3416
rect -5264 -3416 -5194 -2984
rect -5098 2984 -5028 3416
rect -5098 -3416 -5028 -2984
rect -4932 2984 -4862 3416
rect -4932 -3416 -4862 -2984
rect -4766 2984 -4696 3416
rect -4766 -3416 -4696 -2984
rect -4600 2984 -4530 3416
rect -4600 -3416 -4530 -2984
rect -4434 2984 -4364 3416
rect -4434 -3416 -4364 -2984
rect -4268 2984 -4198 3416
rect -4268 -3416 -4198 -2984
rect -4102 2984 -4032 3416
rect -4102 -3416 -4032 -2984
rect -3936 2984 -3866 3416
rect -3936 -3416 -3866 -2984
rect -3770 2984 -3700 3416
rect -3770 -3416 -3700 -2984
rect -3604 2984 -3534 3416
rect -3604 -3416 -3534 -2984
rect -3438 2984 -3368 3416
rect -3438 -3416 -3368 -2984
rect -3272 2984 -3202 3416
rect -3272 -3416 -3202 -2984
rect -3106 2984 -3036 3416
rect -3106 -3416 -3036 -2984
rect -2940 2984 -2870 3416
rect -2940 -3416 -2870 -2984
rect -2774 2984 -2704 3416
rect -2774 -3416 -2704 -2984
rect -2608 2984 -2538 3416
rect -2608 -3416 -2538 -2984
rect -2442 2984 -2372 3416
rect -2442 -3416 -2372 -2984
rect -2276 2984 -2206 3416
rect -2276 -3416 -2206 -2984
rect -2110 2984 -2040 3416
rect -2110 -3416 -2040 -2984
rect -1944 2984 -1874 3416
rect -1944 -3416 -1874 -2984
rect -1778 2984 -1708 3416
rect -1778 -3416 -1708 -2984
rect -1612 2984 -1542 3416
rect -1612 -3416 -1542 -2984
rect -1446 2984 -1376 3416
rect -1446 -3416 -1376 -2984
rect -1280 2984 -1210 3416
rect -1280 -3416 -1210 -2984
rect -1114 2984 -1044 3416
rect -1114 -3416 -1044 -2984
rect -948 2984 -878 3416
rect -948 -3416 -878 -2984
rect -782 2984 -712 3416
rect -782 -3416 -712 -2984
rect -616 2984 -546 3416
rect -616 -3416 -546 -2984
rect -450 2984 -380 3416
rect -450 -3416 -380 -2984
rect -284 2984 -214 3416
rect -284 -3416 -214 -2984
rect -118 2984 -48 3416
rect -118 -3416 -48 -2984
rect 48 2984 118 3416
rect 48 -3416 118 -2984
rect 214 2984 284 3416
rect 214 -3416 284 -2984
rect 380 2984 450 3416
rect 380 -3416 450 -2984
rect 546 2984 616 3416
rect 546 -3416 616 -2984
rect 712 2984 782 3416
rect 712 -3416 782 -2984
rect 878 2984 948 3416
rect 878 -3416 948 -2984
rect 1044 2984 1114 3416
rect 1044 -3416 1114 -2984
rect 1210 2984 1280 3416
rect 1210 -3416 1280 -2984
rect 1376 2984 1446 3416
rect 1376 -3416 1446 -2984
rect 1542 2984 1612 3416
rect 1542 -3416 1612 -2984
rect 1708 2984 1778 3416
rect 1708 -3416 1778 -2984
rect 1874 2984 1944 3416
rect 1874 -3416 1944 -2984
rect 2040 2984 2110 3416
rect 2040 -3416 2110 -2984
rect 2206 2984 2276 3416
rect 2206 -3416 2276 -2984
rect 2372 2984 2442 3416
rect 2372 -3416 2442 -2984
rect 2538 2984 2608 3416
rect 2538 -3416 2608 -2984
rect 2704 2984 2774 3416
rect 2704 -3416 2774 -2984
rect 2870 2984 2940 3416
rect 2870 -3416 2940 -2984
rect 3036 2984 3106 3416
rect 3036 -3416 3106 -2984
rect 3202 2984 3272 3416
rect 3202 -3416 3272 -2984
rect 3368 2984 3438 3416
rect 3368 -3416 3438 -2984
rect 3534 2984 3604 3416
rect 3534 -3416 3604 -2984
rect 3700 2984 3770 3416
rect 3700 -3416 3770 -2984
rect 3866 2984 3936 3416
rect 3866 -3416 3936 -2984
rect 4032 2984 4102 3416
rect 4032 -3416 4102 -2984
rect 4198 2984 4268 3416
rect 4198 -3416 4268 -2984
rect 4364 2984 4434 3416
rect 4364 -3416 4434 -2984
rect 4530 2984 4600 3416
rect 4530 -3416 4600 -2984
rect 4696 2984 4766 3416
rect 4696 -3416 4766 -2984
rect 4862 2984 4932 3416
rect 4862 -3416 4932 -2984
rect 5028 2984 5098 3416
rect 5028 -3416 5098 -2984
rect 5194 2984 5264 3416
rect 5194 -3416 5264 -2984
rect 5360 2984 5430 3416
rect 5360 -3416 5430 -2984
rect 5526 2984 5596 3416
rect 5526 -3416 5596 -2984
rect 5692 2984 5762 3416
rect 5692 -3416 5762 -2984
rect 5858 2984 5928 3416
rect 5858 -3416 5928 -2984
rect 6024 2984 6094 3416
rect 6024 -3416 6094 -2984
rect 6190 2984 6260 3416
rect 6190 -3416 6260 -2984
rect 6356 2984 6426 3416
rect 6356 -3416 6426 -2984
rect 6522 2984 6592 3416
rect 6522 -3416 6592 -2984
<< ppolyres >>
rect -6592 -2984 -6522 2984
rect -6426 -2984 -6356 2984
rect -6260 -2984 -6190 2984
rect -6094 -2984 -6024 2984
rect -5928 -2984 -5858 2984
rect -5762 -2984 -5692 2984
rect -5596 -2984 -5526 2984
rect -5430 -2984 -5360 2984
rect -5264 -2984 -5194 2984
rect -5098 -2984 -5028 2984
rect -4932 -2984 -4862 2984
rect -4766 -2984 -4696 2984
rect -4600 -2984 -4530 2984
rect -4434 -2984 -4364 2984
rect -4268 -2984 -4198 2984
rect -4102 -2984 -4032 2984
rect -3936 -2984 -3866 2984
rect -3770 -2984 -3700 2984
rect -3604 -2984 -3534 2984
rect -3438 -2984 -3368 2984
rect -3272 -2984 -3202 2984
rect -3106 -2984 -3036 2984
rect -2940 -2984 -2870 2984
rect -2774 -2984 -2704 2984
rect -2608 -2984 -2538 2984
rect -2442 -2984 -2372 2984
rect -2276 -2984 -2206 2984
rect -2110 -2984 -2040 2984
rect -1944 -2984 -1874 2984
rect -1778 -2984 -1708 2984
rect -1612 -2984 -1542 2984
rect -1446 -2984 -1376 2984
rect -1280 -2984 -1210 2984
rect -1114 -2984 -1044 2984
rect -948 -2984 -878 2984
rect -782 -2984 -712 2984
rect -616 -2984 -546 2984
rect -450 -2984 -380 2984
rect -284 -2984 -214 2984
rect -118 -2984 -48 2984
rect 48 -2984 118 2984
rect 214 -2984 284 2984
rect 380 -2984 450 2984
rect 546 -2984 616 2984
rect 712 -2984 782 2984
rect 878 -2984 948 2984
rect 1044 -2984 1114 2984
rect 1210 -2984 1280 2984
rect 1376 -2984 1446 2984
rect 1542 -2984 1612 2984
rect 1708 -2984 1778 2984
rect 1874 -2984 1944 2984
rect 2040 -2984 2110 2984
rect 2206 -2984 2276 2984
rect 2372 -2984 2442 2984
rect 2538 -2984 2608 2984
rect 2704 -2984 2774 2984
rect 2870 -2984 2940 2984
rect 3036 -2984 3106 2984
rect 3202 -2984 3272 2984
rect 3368 -2984 3438 2984
rect 3534 -2984 3604 2984
rect 3700 -2984 3770 2984
rect 3866 -2984 3936 2984
rect 4032 -2984 4102 2984
rect 4198 -2984 4268 2984
rect 4364 -2984 4434 2984
rect 4530 -2984 4600 2984
rect 4696 -2984 4766 2984
rect 4862 -2984 4932 2984
rect 5028 -2984 5098 2984
rect 5194 -2984 5264 2984
rect 5360 -2984 5430 2984
rect 5526 -2984 5596 2984
rect 5692 -2984 5762 2984
rect 5858 -2984 5928 2984
rect 6024 -2984 6094 2984
rect 6190 -2984 6260 2984
rect 6356 -2984 6426 2984
rect 6522 -2984 6592 2984
<< locali >>
rect -6722 3512 -6626 3546
rect 6626 3512 6722 3546
rect -6722 3450 -6688 3512
rect 6688 3450 6722 3512
rect -6722 -3512 -6688 -3450
rect 6688 -3512 6722 -3450
rect -6722 -3546 -6626 -3512
rect 6626 -3546 6722 -3512
<< viali >>
rect -6019 3512 6019 3546
rect -6722 -3161 -6688 3161
rect -6576 3001 -6538 3398
rect -6410 3001 -6372 3398
rect -6244 3001 -6206 3398
rect -6078 3001 -6040 3398
rect -5912 3001 -5874 3398
rect -5746 3001 -5708 3398
rect -5580 3001 -5542 3398
rect -5414 3001 -5376 3398
rect -5248 3001 -5210 3398
rect -5082 3001 -5044 3398
rect -4916 3001 -4878 3398
rect -4750 3001 -4712 3398
rect -4584 3001 -4546 3398
rect -4418 3001 -4380 3398
rect -4252 3001 -4214 3398
rect -4086 3001 -4048 3398
rect -3920 3001 -3882 3398
rect -3754 3001 -3716 3398
rect -3588 3001 -3550 3398
rect -3422 3001 -3384 3398
rect -3256 3001 -3218 3398
rect -3090 3001 -3052 3398
rect -2924 3001 -2886 3398
rect -2758 3001 -2720 3398
rect -2592 3001 -2554 3398
rect -2426 3001 -2388 3398
rect -2260 3001 -2222 3398
rect -2094 3001 -2056 3398
rect -1928 3001 -1890 3398
rect -1762 3001 -1724 3398
rect -1596 3001 -1558 3398
rect -1430 3001 -1392 3398
rect -1264 3001 -1226 3398
rect -1098 3001 -1060 3398
rect -932 3001 -894 3398
rect -766 3001 -728 3398
rect -600 3001 -562 3398
rect -434 3001 -396 3398
rect -268 3001 -230 3398
rect -102 3001 -64 3398
rect 64 3001 102 3398
rect 230 3001 268 3398
rect 396 3001 434 3398
rect 562 3001 600 3398
rect 728 3001 766 3398
rect 894 3001 932 3398
rect 1060 3001 1098 3398
rect 1226 3001 1264 3398
rect 1392 3001 1430 3398
rect 1558 3001 1596 3398
rect 1724 3001 1762 3398
rect 1890 3001 1928 3398
rect 2056 3001 2094 3398
rect 2222 3001 2260 3398
rect 2388 3001 2426 3398
rect 2554 3001 2592 3398
rect 2720 3001 2758 3398
rect 2886 3001 2924 3398
rect 3052 3001 3090 3398
rect 3218 3001 3256 3398
rect 3384 3001 3422 3398
rect 3550 3001 3588 3398
rect 3716 3001 3754 3398
rect 3882 3001 3920 3398
rect 4048 3001 4086 3398
rect 4214 3001 4252 3398
rect 4380 3001 4418 3398
rect 4546 3001 4584 3398
rect 4712 3001 4750 3398
rect 4878 3001 4916 3398
rect 5044 3001 5082 3398
rect 5210 3001 5248 3398
rect 5376 3001 5414 3398
rect 5542 3001 5580 3398
rect 5708 3001 5746 3398
rect 5874 3001 5912 3398
rect 6040 3001 6078 3398
rect 6206 3001 6244 3398
rect 6372 3001 6410 3398
rect 6538 3001 6576 3398
rect 6688 -2810 6722 2810
rect -6576 -3398 -6538 -3001
rect -6410 -3398 -6372 -3001
rect -6244 -3398 -6206 -3001
rect -6078 -3398 -6040 -3001
rect -5912 -3398 -5874 -3001
rect -5746 -3398 -5708 -3001
rect -5580 -3398 -5542 -3001
rect -5414 -3398 -5376 -3001
rect -5248 -3398 -5210 -3001
rect -5082 -3398 -5044 -3001
rect -4916 -3398 -4878 -3001
rect -4750 -3398 -4712 -3001
rect -4584 -3398 -4546 -3001
rect -4418 -3398 -4380 -3001
rect -4252 -3398 -4214 -3001
rect -4086 -3398 -4048 -3001
rect -3920 -3398 -3882 -3001
rect -3754 -3398 -3716 -3001
rect -3588 -3398 -3550 -3001
rect -3422 -3398 -3384 -3001
rect -3256 -3398 -3218 -3001
rect -3090 -3398 -3052 -3001
rect -2924 -3398 -2886 -3001
rect -2758 -3398 -2720 -3001
rect -2592 -3398 -2554 -3001
rect -2426 -3398 -2388 -3001
rect -2260 -3398 -2222 -3001
rect -2094 -3398 -2056 -3001
rect -1928 -3398 -1890 -3001
rect -1762 -3398 -1724 -3001
rect -1596 -3398 -1558 -3001
rect -1430 -3398 -1392 -3001
rect -1264 -3398 -1226 -3001
rect -1098 -3398 -1060 -3001
rect -932 -3398 -894 -3001
rect -766 -3398 -728 -3001
rect -600 -3398 -562 -3001
rect -434 -3398 -396 -3001
rect -268 -3398 -230 -3001
rect -102 -3398 -64 -3001
rect 64 -3398 102 -3001
rect 230 -3398 268 -3001
rect 396 -3398 434 -3001
rect 562 -3398 600 -3001
rect 728 -3398 766 -3001
rect 894 -3398 932 -3001
rect 1060 -3398 1098 -3001
rect 1226 -3398 1264 -3001
rect 1392 -3398 1430 -3001
rect 1558 -3398 1596 -3001
rect 1724 -3398 1762 -3001
rect 1890 -3398 1928 -3001
rect 2056 -3398 2094 -3001
rect 2222 -3398 2260 -3001
rect 2388 -3398 2426 -3001
rect 2554 -3398 2592 -3001
rect 2720 -3398 2758 -3001
rect 2886 -3398 2924 -3001
rect 3052 -3398 3090 -3001
rect 3218 -3398 3256 -3001
rect 3384 -3398 3422 -3001
rect 3550 -3398 3588 -3001
rect 3716 -3398 3754 -3001
rect 3882 -3398 3920 -3001
rect 4048 -3398 4086 -3001
rect 4214 -3398 4252 -3001
rect 4380 -3398 4418 -3001
rect 4546 -3398 4584 -3001
rect 4712 -3398 4750 -3001
rect 4878 -3398 4916 -3001
rect 5044 -3398 5082 -3001
rect 5210 -3398 5248 -3001
rect 5376 -3398 5414 -3001
rect 5542 -3398 5580 -3001
rect 5708 -3398 5746 -3001
rect 5874 -3398 5912 -3001
rect 6040 -3398 6078 -3001
rect 6206 -3398 6244 -3001
rect 6372 -3398 6410 -3001
rect 6538 -3398 6576 -3001
rect -6019 -3546 6019 -3512
<< metal1 >>
rect -6031 3546 6031 3552
rect -6031 3512 -6019 3546
rect 6019 3512 6031 3546
rect -6031 3506 6031 3512
rect -6582 3398 -6532 3410
rect -6728 3161 -6682 3173
rect -6728 -3161 -6722 3161
rect -6688 -3161 -6682 3161
rect -6582 3001 -6576 3398
rect -6538 3001 -6532 3398
rect -6582 2989 -6532 3001
rect -6416 3398 -6366 3410
rect -6416 3001 -6410 3398
rect -6372 3001 -6366 3398
rect -6416 2989 -6366 3001
rect -6250 3398 -6200 3410
rect -6250 3001 -6244 3398
rect -6206 3001 -6200 3398
rect -6250 2989 -6200 3001
rect -6084 3398 -6034 3410
rect -6084 3001 -6078 3398
rect -6040 3001 -6034 3398
rect -6084 2989 -6034 3001
rect -5918 3398 -5868 3410
rect -5918 3001 -5912 3398
rect -5874 3001 -5868 3398
rect -5918 2989 -5868 3001
rect -5752 3398 -5702 3410
rect -5752 3001 -5746 3398
rect -5708 3001 -5702 3398
rect -5752 2989 -5702 3001
rect -5586 3398 -5536 3410
rect -5586 3001 -5580 3398
rect -5542 3001 -5536 3398
rect -5586 2989 -5536 3001
rect -5420 3398 -5370 3410
rect -5420 3001 -5414 3398
rect -5376 3001 -5370 3398
rect -5420 2989 -5370 3001
rect -5254 3398 -5204 3410
rect -5254 3001 -5248 3398
rect -5210 3001 -5204 3398
rect -5254 2989 -5204 3001
rect -5088 3398 -5038 3410
rect -5088 3001 -5082 3398
rect -5044 3001 -5038 3398
rect -5088 2989 -5038 3001
rect -4922 3398 -4872 3410
rect -4922 3001 -4916 3398
rect -4878 3001 -4872 3398
rect -4922 2989 -4872 3001
rect -4756 3398 -4706 3410
rect -4756 3001 -4750 3398
rect -4712 3001 -4706 3398
rect -4756 2989 -4706 3001
rect -4590 3398 -4540 3410
rect -4590 3001 -4584 3398
rect -4546 3001 -4540 3398
rect -4590 2989 -4540 3001
rect -4424 3398 -4374 3410
rect -4424 3001 -4418 3398
rect -4380 3001 -4374 3398
rect -4424 2989 -4374 3001
rect -4258 3398 -4208 3410
rect -4258 3001 -4252 3398
rect -4214 3001 -4208 3398
rect -4258 2989 -4208 3001
rect -4092 3398 -4042 3410
rect -4092 3001 -4086 3398
rect -4048 3001 -4042 3398
rect -4092 2989 -4042 3001
rect -3926 3398 -3876 3410
rect -3926 3001 -3920 3398
rect -3882 3001 -3876 3398
rect -3926 2989 -3876 3001
rect -3760 3398 -3710 3410
rect -3760 3001 -3754 3398
rect -3716 3001 -3710 3398
rect -3760 2989 -3710 3001
rect -3594 3398 -3544 3410
rect -3594 3001 -3588 3398
rect -3550 3001 -3544 3398
rect -3594 2989 -3544 3001
rect -3428 3398 -3378 3410
rect -3428 3001 -3422 3398
rect -3384 3001 -3378 3398
rect -3428 2989 -3378 3001
rect -3262 3398 -3212 3410
rect -3262 3001 -3256 3398
rect -3218 3001 -3212 3398
rect -3262 2989 -3212 3001
rect -3096 3398 -3046 3410
rect -3096 3001 -3090 3398
rect -3052 3001 -3046 3398
rect -3096 2989 -3046 3001
rect -2930 3398 -2880 3410
rect -2930 3001 -2924 3398
rect -2886 3001 -2880 3398
rect -2930 2989 -2880 3001
rect -2764 3398 -2714 3410
rect -2764 3001 -2758 3398
rect -2720 3001 -2714 3398
rect -2764 2989 -2714 3001
rect -2598 3398 -2548 3410
rect -2598 3001 -2592 3398
rect -2554 3001 -2548 3398
rect -2598 2989 -2548 3001
rect -2432 3398 -2382 3410
rect -2432 3001 -2426 3398
rect -2388 3001 -2382 3398
rect -2432 2989 -2382 3001
rect -2266 3398 -2216 3410
rect -2266 3001 -2260 3398
rect -2222 3001 -2216 3398
rect -2266 2989 -2216 3001
rect -2100 3398 -2050 3410
rect -2100 3001 -2094 3398
rect -2056 3001 -2050 3398
rect -2100 2989 -2050 3001
rect -1934 3398 -1884 3410
rect -1934 3001 -1928 3398
rect -1890 3001 -1884 3398
rect -1934 2989 -1884 3001
rect -1768 3398 -1718 3410
rect -1768 3001 -1762 3398
rect -1724 3001 -1718 3398
rect -1768 2989 -1718 3001
rect -1602 3398 -1552 3410
rect -1602 3001 -1596 3398
rect -1558 3001 -1552 3398
rect -1602 2989 -1552 3001
rect -1436 3398 -1386 3410
rect -1436 3001 -1430 3398
rect -1392 3001 -1386 3398
rect -1436 2989 -1386 3001
rect -1270 3398 -1220 3410
rect -1270 3001 -1264 3398
rect -1226 3001 -1220 3398
rect -1270 2989 -1220 3001
rect -1104 3398 -1054 3410
rect -1104 3001 -1098 3398
rect -1060 3001 -1054 3398
rect -1104 2989 -1054 3001
rect -938 3398 -888 3410
rect -938 3001 -932 3398
rect -894 3001 -888 3398
rect -938 2989 -888 3001
rect -772 3398 -722 3410
rect -772 3001 -766 3398
rect -728 3001 -722 3398
rect -772 2989 -722 3001
rect -606 3398 -556 3410
rect -606 3001 -600 3398
rect -562 3001 -556 3398
rect -606 2989 -556 3001
rect -440 3398 -390 3410
rect -440 3001 -434 3398
rect -396 3001 -390 3398
rect -440 2989 -390 3001
rect -274 3398 -224 3410
rect -274 3001 -268 3398
rect -230 3001 -224 3398
rect -274 2989 -224 3001
rect -108 3398 -58 3410
rect -108 3001 -102 3398
rect -64 3001 -58 3398
rect -108 2989 -58 3001
rect 58 3398 108 3410
rect 58 3001 64 3398
rect 102 3001 108 3398
rect 58 2989 108 3001
rect 224 3398 274 3410
rect 224 3001 230 3398
rect 268 3001 274 3398
rect 224 2989 274 3001
rect 390 3398 440 3410
rect 390 3001 396 3398
rect 434 3001 440 3398
rect 390 2989 440 3001
rect 556 3398 606 3410
rect 556 3001 562 3398
rect 600 3001 606 3398
rect 556 2989 606 3001
rect 722 3398 772 3410
rect 722 3001 728 3398
rect 766 3001 772 3398
rect 722 2989 772 3001
rect 888 3398 938 3410
rect 888 3001 894 3398
rect 932 3001 938 3398
rect 888 2989 938 3001
rect 1054 3398 1104 3410
rect 1054 3001 1060 3398
rect 1098 3001 1104 3398
rect 1054 2989 1104 3001
rect 1220 3398 1270 3410
rect 1220 3001 1226 3398
rect 1264 3001 1270 3398
rect 1220 2989 1270 3001
rect 1386 3398 1436 3410
rect 1386 3001 1392 3398
rect 1430 3001 1436 3398
rect 1386 2989 1436 3001
rect 1552 3398 1602 3410
rect 1552 3001 1558 3398
rect 1596 3001 1602 3398
rect 1552 2989 1602 3001
rect 1718 3398 1768 3410
rect 1718 3001 1724 3398
rect 1762 3001 1768 3398
rect 1718 2989 1768 3001
rect 1884 3398 1934 3410
rect 1884 3001 1890 3398
rect 1928 3001 1934 3398
rect 1884 2989 1934 3001
rect 2050 3398 2100 3410
rect 2050 3001 2056 3398
rect 2094 3001 2100 3398
rect 2050 2989 2100 3001
rect 2216 3398 2266 3410
rect 2216 3001 2222 3398
rect 2260 3001 2266 3398
rect 2216 2989 2266 3001
rect 2382 3398 2432 3410
rect 2382 3001 2388 3398
rect 2426 3001 2432 3398
rect 2382 2989 2432 3001
rect 2548 3398 2598 3410
rect 2548 3001 2554 3398
rect 2592 3001 2598 3398
rect 2548 2989 2598 3001
rect 2714 3398 2764 3410
rect 2714 3001 2720 3398
rect 2758 3001 2764 3398
rect 2714 2989 2764 3001
rect 2880 3398 2930 3410
rect 2880 3001 2886 3398
rect 2924 3001 2930 3398
rect 2880 2989 2930 3001
rect 3046 3398 3096 3410
rect 3046 3001 3052 3398
rect 3090 3001 3096 3398
rect 3046 2989 3096 3001
rect 3212 3398 3262 3410
rect 3212 3001 3218 3398
rect 3256 3001 3262 3398
rect 3212 2989 3262 3001
rect 3378 3398 3428 3410
rect 3378 3001 3384 3398
rect 3422 3001 3428 3398
rect 3378 2989 3428 3001
rect 3544 3398 3594 3410
rect 3544 3001 3550 3398
rect 3588 3001 3594 3398
rect 3544 2989 3594 3001
rect 3710 3398 3760 3410
rect 3710 3001 3716 3398
rect 3754 3001 3760 3398
rect 3710 2989 3760 3001
rect 3876 3398 3926 3410
rect 3876 3001 3882 3398
rect 3920 3001 3926 3398
rect 3876 2989 3926 3001
rect 4042 3398 4092 3410
rect 4042 3001 4048 3398
rect 4086 3001 4092 3398
rect 4042 2989 4092 3001
rect 4208 3398 4258 3410
rect 4208 3001 4214 3398
rect 4252 3001 4258 3398
rect 4208 2989 4258 3001
rect 4374 3398 4424 3410
rect 4374 3001 4380 3398
rect 4418 3001 4424 3398
rect 4374 2989 4424 3001
rect 4540 3398 4590 3410
rect 4540 3001 4546 3398
rect 4584 3001 4590 3398
rect 4540 2989 4590 3001
rect 4706 3398 4756 3410
rect 4706 3001 4712 3398
rect 4750 3001 4756 3398
rect 4706 2989 4756 3001
rect 4872 3398 4922 3410
rect 4872 3001 4878 3398
rect 4916 3001 4922 3398
rect 4872 2989 4922 3001
rect 5038 3398 5088 3410
rect 5038 3001 5044 3398
rect 5082 3001 5088 3398
rect 5038 2989 5088 3001
rect 5204 3398 5254 3410
rect 5204 3001 5210 3398
rect 5248 3001 5254 3398
rect 5204 2989 5254 3001
rect 5370 3398 5420 3410
rect 5370 3001 5376 3398
rect 5414 3001 5420 3398
rect 5370 2989 5420 3001
rect 5536 3398 5586 3410
rect 5536 3001 5542 3398
rect 5580 3001 5586 3398
rect 5536 2989 5586 3001
rect 5702 3398 5752 3410
rect 5702 3001 5708 3398
rect 5746 3001 5752 3398
rect 5702 2989 5752 3001
rect 5868 3398 5918 3410
rect 5868 3001 5874 3398
rect 5912 3001 5918 3398
rect 5868 2989 5918 3001
rect 6034 3398 6084 3410
rect 6034 3001 6040 3398
rect 6078 3001 6084 3398
rect 6034 2989 6084 3001
rect 6200 3398 6250 3410
rect 6200 3001 6206 3398
rect 6244 3001 6250 3398
rect 6200 2989 6250 3001
rect 6366 3398 6416 3410
rect 6366 3001 6372 3398
rect 6410 3001 6416 3398
rect 6366 2989 6416 3001
rect 6532 3398 6582 3410
rect 6532 3001 6538 3398
rect 6576 3001 6582 3398
rect 6532 2989 6582 3001
rect 6682 2810 6728 2822
rect 6682 -2810 6688 2810
rect 6722 -2810 6728 2810
rect 6682 -2822 6728 -2810
rect -6728 -3173 -6682 -3161
rect -6582 -3001 -6532 -2989
rect -6582 -3398 -6576 -3001
rect -6538 -3398 -6532 -3001
rect -6582 -3410 -6532 -3398
rect -6416 -3001 -6366 -2989
rect -6416 -3398 -6410 -3001
rect -6372 -3398 -6366 -3001
rect -6416 -3410 -6366 -3398
rect -6250 -3001 -6200 -2989
rect -6250 -3398 -6244 -3001
rect -6206 -3398 -6200 -3001
rect -6250 -3410 -6200 -3398
rect -6084 -3001 -6034 -2989
rect -6084 -3398 -6078 -3001
rect -6040 -3398 -6034 -3001
rect -6084 -3410 -6034 -3398
rect -5918 -3001 -5868 -2989
rect -5918 -3398 -5912 -3001
rect -5874 -3398 -5868 -3001
rect -5918 -3410 -5868 -3398
rect -5752 -3001 -5702 -2989
rect -5752 -3398 -5746 -3001
rect -5708 -3398 -5702 -3001
rect -5752 -3410 -5702 -3398
rect -5586 -3001 -5536 -2989
rect -5586 -3398 -5580 -3001
rect -5542 -3398 -5536 -3001
rect -5586 -3410 -5536 -3398
rect -5420 -3001 -5370 -2989
rect -5420 -3398 -5414 -3001
rect -5376 -3398 -5370 -3001
rect -5420 -3410 -5370 -3398
rect -5254 -3001 -5204 -2989
rect -5254 -3398 -5248 -3001
rect -5210 -3398 -5204 -3001
rect -5254 -3410 -5204 -3398
rect -5088 -3001 -5038 -2989
rect -5088 -3398 -5082 -3001
rect -5044 -3398 -5038 -3001
rect -5088 -3410 -5038 -3398
rect -4922 -3001 -4872 -2989
rect -4922 -3398 -4916 -3001
rect -4878 -3398 -4872 -3001
rect -4922 -3410 -4872 -3398
rect -4756 -3001 -4706 -2989
rect -4756 -3398 -4750 -3001
rect -4712 -3398 -4706 -3001
rect -4756 -3410 -4706 -3398
rect -4590 -3001 -4540 -2989
rect -4590 -3398 -4584 -3001
rect -4546 -3398 -4540 -3001
rect -4590 -3410 -4540 -3398
rect -4424 -3001 -4374 -2989
rect -4424 -3398 -4418 -3001
rect -4380 -3398 -4374 -3001
rect -4424 -3410 -4374 -3398
rect -4258 -3001 -4208 -2989
rect -4258 -3398 -4252 -3001
rect -4214 -3398 -4208 -3001
rect -4258 -3410 -4208 -3398
rect -4092 -3001 -4042 -2989
rect -4092 -3398 -4086 -3001
rect -4048 -3398 -4042 -3001
rect -4092 -3410 -4042 -3398
rect -3926 -3001 -3876 -2989
rect -3926 -3398 -3920 -3001
rect -3882 -3398 -3876 -3001
rect -3926 -3410 -3876 -3398
rect -3760 -3001 -3710 -2989
rect -3760 -3398 -3754 -3001
rect -3716 -3398 -3710 -3001
rect -3760 -3410 -3710 -3398
rect -3594 -3001 -3544 -2989
rect -3594 -3398 -3588 -3001
rect -3550 -3398 -3544 -3001
rect -3594 -3410 -3544 -3398
rect -3428 -3001 -3378 -2989
rect -3428 -3398 -3422 -3001
rect -3384 -3398 -3378 -3001
rect -3428 -3410 -3378 -3398
rect -3262 -3001 -3212 -2989
rect -3262 -3398 -3256 -3001
rect -3218 -3398 -3212 -3001
rect -3262 -3410 -3212 -3398
rect -3096 -3001 -3046 -2989
rect -3096 -3398 -3090 -3001
rect -3052 -3398 -3046 -3001
rect -3096 -3410 -3046 -3398
rect -2930 -3001 -2880 -2989
rect -2930 -3398 -2924 -3001
rect -2886 -3398 -2880 -3001
rect -2930 -3410 -2880 -3398
rect -2764 -3001 -2714 -2989
rect -2764 -3398 -2758 -3001
rect -2720 -3398 -2714 -3001
rect -2764 -3410 -2714 -3398
rect -2598 -3001 -2548 -2989
rect -2598 -3398 -2592 -3001
rect -2554 -3398 -2548 -3001
rect -2598 -3410 -2548 -3398
rect -2432 -3001 -2382 -2989
rect -2432 -3398 -2426 -3001
rect -2388 -3398 -2382 -3001
rect -2432 -3410 -2382 -3398
rect -2266 -3001 -2216 -2989
rect -2266 -3398 -2260 -3001
rect -2222 -3398 -2216 -3001
rect -2266 -3410 -2216 -3398
rect -2100 -3001 -2050 -2989
rect -2100 -3398 -2094 -3001
rect -2056 -3398 -2050 -3001
rect -2100 -3410 -2050 -3398
rect -1934 -3001 -1884 -2989
rect -1934 -3398 -1928 -3001
rect -1890 -3398 -1884 -3001
rect -1934 -3410 -1884 -3398
rect -1768 -3001 -1718 -2989
rect -1768 -3398 -1762 -3001
rect -1724 -3398 -1718 -3001
rect -1768 -3410 -1718 -3398
rect -1602 -3001 -1552 -2989
rect -1602 -3398 -1596 -3001
rect -1558 -3398 -1552 -3001
rect -1602 -3410 -1552 -3398
rect -1436 -3001 -1386 -2989
rect -1436 -3398 -1430 -3001
rect -1392 -3398 -1386 -3001
rect -1436 -3410 -1386 -3398
rect -1270 -3001 -1220 -2989
rect -1270 -3398 -1264 -3001
rect -1226 -3398 -1220 -3001
rect -1270 -3410 -1220 -3398
rect -1104 -3001 -1054 -2989
rect -1104 -3398 -1098 -3001
rect -1060 -3398 -1054 -3001
rect -1104 -3410 -1054 -3398
rect -938 -3001 -888 -2989
rect -938 -3398 -932 -3001
rect -894 -3398 -888 -3001
rect -938 -3410 -888 -3398
rect -772 -3001 -722 -2989
rect -772 -3398 -766 -3001
rect -728 -3398 -722 -3001
rect -772 -3410 -722 -3398
rect -606 -3001 -556 -2989
rect -606 -3398 -600 -3001
rect -562 -3398 -556 -3001
rect -606 -3410 -556 -3398
rect -440 -3001 -390 -2989
rect -440 -3398 -434 -3001
rect -396 -3398 -390 -3001
rect -440 -3410 -390 -3398
rect -274 -3001 -224 -2989
rect -274 -3398 -268 -3001
rect -230 -3398 -224 -3001
rect -274 -3410 -224 -3398
rect -108 -3001 -58 -2989
rect -108 -3398 -102 -3001
rect -64 -3398 -58 -3001
rect -108 -3410 -58 -3398
rect 58 -3001 108 -2989
rect 58 -3398 64 -3001
rect 102 -3398 108 -3001
rect 58 -3410 108 -3398
rect 224 -3001 274 -2989
rect 224 -3398 230 -3001
rect 268 -3398 274 -3001
rect 224 -3410 274 -3398
rect 390 -3001 440 -2989
rect 390 -3398 396 -3001
rect 434 -3398 440 -3001
rect 390 -3410 440 -3398
rect 556 -3001 606 -2989
rect 556 -3398 562 -3001
rect 600 -3398 606 -3001
rect 556 -3410 606 -3398
rect 722 -3001 772 -2989
rect 722 -3398 728 -3001
rect 766 -3398 772 -3001
rect 722 -3410 772 -3398
rect 888 -3001 938 -2989
rect 888 -3398 894 -3001
rect 932 -3398 938 -3001
rect 888 -3410 938 -3398
rect 1054 -3001 1104 -2989
rect 1054 -3398 1060 -3001
rect 1098 -3398 1104 -3001
rect 1054 -3410 1104 -3398
rect 1220 -3001 1270 -2989
rect 1220 -3398 1226 -3001
rect 1264 -3398 1270 -3001
rect 1220 -3410 1270 -3398
rect 1386 -3001 1436 -2989
rect 1386 -3398 1392 -3001
rect 1430 -3398 1436 -3001
rect 1386 -3410 1436 -3398
rect 1552 -3001 1602 -2989
rect 1552 -3398 1558 -3001
rect 1596 -3398 1602 -3001
rect 1552 -3410 1602 -3398
rect 1718 -3001 1768 -2989
rect 1718 -3398 1724 -3001
rect 1762 -3398 1768 -3001
rect 1718 -3410 1768 -3398
rect 1884 -3001 1934 -2989
rect 1884 -3398 1890 -3001
rect 1928 -3398 1934 -3001
rect 1884 -3410 1934 -3398
rect 2050 -3001 2100 -2989
rect 2050 -3398 2056 -3001
rect 2094 -3398 2100 -3001
rect 2050 -3410 2100 -3398
rect 2216 -3001 2266 -2989
rect 2216 -3398 2222 -3001
rect 2260 -3398 2266 -3001
rect 2216 -3410 2266 -3398
rect 2382 -3001 2432 -2989
rect 2382 -3398 2388 -3001
rect 2426 -3398 2432 -3001
rect 2382 -3410 2432 -3398
rect 2548 -3001 2598 -2989
rect 2548 -3398 2554 -3001
rect 2592 -3398 2598 -3001
rect 2548 -3410 2598 -3398
rect 2714 -3001 2764 -2989
rect 2714 -3398 2720 -3001
rect 2758 -3398 2764 -3001
rect 2714 -3410 2764 -3398
rect 2880 -3001 2930 -2989
rect 2880 -3398 2886 -3001
rect 2924 -3398 2930 -3001
rect 2880 -3410 2930 -3398
rect 3046 -3001 3096 -2989
rect 3046 -3398 3052 -3001
rect 3090 -3398 3096 -3001
rect 3046 -3410 3096 -3398
rect 3212 -3001 3262 -2989
rect 3212 -3398 3218 -3001
rect 3256 -3398 3262 -3001
rect 3212 -3410 3262 -3398
rect 3378 -3001 3428 -2989
rect 3378 -3398 3384 -3001
rect 3422 -3398 3428 -3001
rect 3378 -3410 3428 -3398
rect 3544 -3001 3594 -2989
rect 3544 -3398 3550 -3001
rect 3588 -3398 3594 -3001
rect 3544 -3410 3594 -3398
rect 3710 -3001 3760 -2989
rect 3710 -3398 3716 -3001
rect 3754 -3398 3760 -3001
rect 3710 -3410 3760 -3398
rect 3876 -3001 3926 -2989
rect 3876 -3398 3882 -3001
rect 3920 -3398 3926 -3001
rect 3876 -3410 3926 -3398
rect 4042 -3001 4092 -2989
rect 4042 -3398 4048 -3001
rect 4086 -3398 4092 -3001
rect 4042 -3410 4092 -3398
rect 4208 -3001 4258 -2989
rect 4208 -3398 4214 -3001
rect 4252 -3398 4258 -3001
rect 4208 -3410 4258 -3398
rect 4374 -3001 4424 -2989
rect 4374 -3398 4380 -3001
rect 4418 -3398 4424 -3001
rect 4374 -3410 4424 -3398
rect 4540 -3001 4590 -2989
rect 4540 -3398 4546 -3001
rect 4584 -3398 4590 -3001
rect 4540 -3410 4590 -3398
rect 4706 -3001 4756 -2989
rect 4706 -3398 4712 -3001
rect 4750 -3398 4756 -3001
rect 4706 -3410 4756 -3398
rect 4872 -3001 4922 -2989
rect 4872 -3398 4878 -3001
rect 4916 -3398 4922 -3001
rect 4872 -3410 4922 -3398
rect 5038 -3001 5088 -2989
rect 5038 -3398 5044 -3001
rect 5082 -3398 5088 -3001
rect 5038 -3410 5088 -3398
rect 5204 -3001 5254 -2989
rect 5204 -3398 5210 -3001
rect 5248 -3398 5254 -3001
rect 5204 -3410 5254 -3398
rect 5370 -3001 5420 -2989
rect 5370 -3398 5376 -3001
rect 5414 -3398 5420 -3001
rect 5370 -3410 5420 -3398
rect 5536 -3001 5586 -2989
rect 5536 -3398 5542 -3001
rect 5580 -3398 5586 -3001
rect 5536 -3410 5586 -3398
rect 5702 -3001 5752 -2989
rect 5702 -3398 5708 -3001
rect 5746 -3398 5752 -3001
rect 5702 -3410 5752 -3398
rect 5868 -3001 5918 -2989
rect 5868 -3398 5874 -3001
rect 5912 -3398 5918 -3001
rect 5868 -3410 5918 -3398
rect 6034 -3001 6084 -2989
rect 6034 -3398 6040 -3001
rect 6078 -3398 6084 -3001
rect 6034 -3410 6084 -3398
rect 6200 -3001 6250 -2989
rect 6200 -3398 6206 -3001
rect 6244 -3398 6250 -3001
rect 6200 -3410 6250 -3398
rect 6366 -3001 6416 -2989
rect 6366 -3398 6372 -3001
rect 6410 -3398 6416 -3001
rect 6366 -3410 6416 -3398
rect 6532 -3001 6582 -2989
rect 6532 -3398 6538 -3001
rect 6576 -3398 6582 -3001
rect 6532 -3410 6582 -3398
rect -6031 -3512 6031 -3506
rect -6031 -3546 -6019 -3512
rect 6019 -3546 6031 -3512
rect -6031 -3552 6031 -3546
<< properties >>
string FIXED_BBOX -6705 -3529 6705 3529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 30.0 m 1 nx 80 wmin 0.350 lmin 0.50 rho 319.8 val 28.524k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 90 viagt 90 viagl 90 viagr 80
<< end >>
