magic
tech sky130A
magscale 1 2
timestamp 1713926953
<< locali >>
rect 3396 364 3448 658
rect 3742 364 3922 658
rect 3396 342 3922 364
rect 3448 270 3742 342
<< metal1 >>
rect 3724 1027 3788 1035
rect 3568 771 3622 777
rect 3304 280 3356 290
rect 3356 144 3357 276
rect 3304 138 3357 144
rect 3305 -1916 3357 138
rect 3392 -1514 3456 52
rect 3568 -610 3622 583
rect 3724 -540 3788 839
rect 3830 282 3882 290
rect 3830 280 3883 282
rect 3882 144 3883 280
rect 3830 138 3883 144
rect 3568 -1622 3620 -860
rect 3305 -2632 3456 -1916
rect 3568 -2584 3620 -1818
rect 3726 -2502 3790 -936
rect 3568 -2586 3616 -2584
rect 3831 -2632 3883 138
rect 3305 -2690 3883 -2632
rect 3304 -2704 3886 -2690
rect 3304 -2782 3362 -2704
rect 3828 -2782 3886 -2704
rect 3304 -2796 3886 -2782
<< via1 >>
rect 3724 839 3788 1027
rect 3568 583 3622 771
rect 3304 144 3356 280
rect 3830 144 3882 280
rect 3568 -1818 3620 -1622
rect 3362 -2782 3828 -2704
<< metal2 >>
rect 3718 839 3724 1027
rect 3788 839 3794 1027
rect 3560 583 3568 771
rect 3622 583 3631 771
rect 3262 280 3922 374
rect 3262 144 3304 280
rect 3356 144 3830 280
rect 3882 144 3922 280
rect 3262 136 3922 144
rect 3262 -852 3922 -614
rect 3262 -1622 3922 -1598
rect 3262 -1818 3568 -1622
rect 3620 -1818 3922 -1622
rect 3262 -1836 3922 -1818
rect 3262 -2704 3922 -2622
rect 3262 -2782 3362 -2704
rect 3828 -2782 3922 -2704
rect 3262 -2860 3922 -2782
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ#1  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 ../../chipalooza/sky130_od_ip__tempsensor/mag
timestamp 1713474431
transform 1 0 3595 0 1 511
box -183 -183 183 183
use sky130_fd_pr__nfet_05v0_nvt_QRKT8P  XM6
timestamp 1713888873
transform 1 0 3594 0 1 -1226
box -328 -558 328 558
use sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P  XM7
timestamp 1713888873
transform 1 0 3594 0 1 -240
box -328 -558 328 558
use sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ  XM12
timestamp 1713896310
transform 1 0 3594 0 1 -2212
box -328 -558 328 558
<< end >>
