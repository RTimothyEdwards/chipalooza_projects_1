magic
tech sky130A
magscale 1 2
timestamp 1713919406
<< error_p >>
rect 561701 354694 561735 354720
rect 561675 354627 561701 354694
rect 561734 354627 561735 354694
rect 561701 354553 561735 354627
rect 561675 353164 561701 354553
rect 561734 353164 561735 354553
rect 561701 349756 561735 350770
rect 561922 349949 561935 350425
rect 561956 349983 561969 350391
rect 561718 349680 561735 349756
rect 561716 348272 561735 349224
rect 561770 348326 561789 349170
rect 561928 348952 561935 349054
rect 561962 348986 561969 349020
rect 561928 348442 561935 348544
rect 561962 348476 561969 348510
rect 561701 348014 561735 348040
rect 561675 347825 561701 348014
rect 561734 347825 561735 348014
rect 561701 347751 561735 347825
rect 561675 347684 561701 347751
rect 561734 347684 561735 347751
rect 561701 345934 561735 345960
rect 561675 345897 561701 345934
rect 561734 345897 561735 345934
rect 561701 345837 561735 345897
rect 562111 345435 565193 345461
rect 565267 345435 565304 345461
rect 562111 345402 562137 345435
rect 562464 345402 562922 345406
rect 564134 345402 564592 345406
rect 565193 345402 565267 345435
rect 562111 345401 565304 345402
rect 565101 344147 565193 344173
rect 565267 344147 565304 344173
rect 565101 344114 565127 344147
rect 565193 344114 565267 344147
rect 565101 344113 565304 344114
rect 564665 343711 564751 343737
rect 564665 343070 564691 343711
rect 564724 343070 564725 343711
rect 564691 341960 564725 341986
rect 564665 341785 564691 341960
rect 564724 341785 564725 341960
rect 564691 341711 564725 341785
rect 564665 341674 564691 341711
rect 564724 341674 564725 341711
rect 51977 254884 52031 254885
rect 51657 254824 51741 254825
rect 51927 254824 51977 254825
rect 56913 49306 56967 49307
rect 56593 49246 56677 49247
rect 56863 49246 56913 49247
rect 273039 10070 273048 10074
rect 273045 10062 273048 10065
rect 273050 10056 273057 10065
rect 273050 10009 273057 10018
rect 273039 10000 273048 10004
rect 138464 1280 138479 1307
rect 138528 1280 138540 1307
rect 141976 1280 141992 1307
rect 145545 1280 145547 1307
rect 149086 1280 149102 1307
rect 152690 1280 152703 1307
rect 188081 1280 188165 1307
rect 191626 1280 191710 1307
rect 195181 1280 195268 1307
rect 138436 1252 138479 1279
rect 138528 1252 138548 1279
rect 141982 1252 141992 1279
rect 145528 1252 145547 1279
rect 149074 1252 149102 1279
rect 152690 1252 152731 1279
rect 188080 1252 188192 1279
rect 191626 1252 191738 1279
rect 195172 1252 195284 1279
rect 191613 983 191626 1010
<< error_s >>
rect 6596 356260 6600 356288
<< metal1 >>
rect 513415 609778 520733 610315
rect 513415 593259 513911 609778
rect 520276 594202 520733 609778
rect 556287 601770 560183 602040
rect 520276 593259 521512 594202
rect 556287 593934 556508 601770
rect 560007 593934 560183 601770
rect 556287 593698 560183 593934
rect 513415 592789 521512 593259
rect 510422 576926 518844 577547
rect 510422 570179 510907 576926
rect 518330 574012 518844 576926
rect 518330 572711 521727 574012
rect 556374 572886 560268 573078
rect 518330 570179 518844 572711
rect 510422 569612 518844 570179
rect 556374 563187 556611 572886
rect 560065 563187 560268 572886
rect 556374 562979 560268 563187
rect 4613 475393 6213 482370
rect 20479 480490 20752 482778
rect 20445 480450 20812 480490
rect 20445 479565 20480 480450
rect 20783 479565 20812 480450
rect 20445 479522 20812 479565
rect 21251 476758 21407 482669
rect 22022 481278 22295 482788
rect 21973 481235 22340 481278
rect 21973 480350 22005 481235
rect 22308 480350 22340 481235
rect 21973 480310 22340 480350
rect 21251 476743 21774 476758
rect 21251 476599 21268 476743
rect 21751 476599 21774 476743
rect 21251 476583 21774 476599
rect 4613 470506 4728 475393
rect 6108 470506 6213 475393
rect 4613 470387 6213 470506
rect 18828 475286 24285 475543
rect 18828 470495 19136 475286
rect 24029 470495 24285 475286
rect 4745 470220 6027 470387
rect 18828 470214 24285 470495
rect 7456 468312 7723 468354
rect 7456 467721 7486 468312
rect 7690 467721 7723 468312
rect 7456 467681 7723 467721
rect 7468 466529 7714 467681
rect 7466 461984 8347 462028
rect 2167 461516 5322 461778
rect 7466 461352 7523 461984
rect 8290 461352 8347 461984
rect 7466 461302 8347 461352
rect 7483 455643 7697 456871
rect 7345 455429 7697 455643
rect 7345 443441 7559 455429
rect 18854 451460 20136 470214
rect 9023 450178 20136 451460
rect 9023 444149 10305 450178
rect 7345 443227 9245 443441
rect 6462 439485 6743 439503
rect 6462 438897 6476 439485
rect 6728 439467 6743 439485
rect 6728 439345 9627 439467
rect 6728 438897 6743 439345
rect 6462 438880 6743 438897
rect 7368 439022 7592 439029
rect 7368 439002 9597 439022
rect 7368 438204 7391 439002
rect 7570 438909 9597 439002
rect 7570 438204 7592 438909
rect 7368 438178 7592 438204
rect 7959 438229 9673 438469
rect 1703 435904 2427 435927
rect 1703 435716 1738 435904
rect 2398 435716 2427 435904
rect 1703 435690 2427 435716
rect 1747 429872 1993 435690
rect 7959 435555 8199 438229
rect 13208 437642 14598 437666
rect 13208 437442 13238 437642
rect 14564 437442 14598 437642
rect 13208 437416 14598 437442
rect 7959 435315 11729 435555
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 6302 429814 7162 429877
rect 11489 429872 11729 435315
rect 4484 426541 4759 426576
rect 4484 425868 4522 426541
rect 4717 426147 4759 426541
rect 6577 426147 6839 427726
rect 4717 425885 6839 426147
rect 4717 425868 4759 425885
rect 4484 425830 4759 425868
rect 580981 367266 581227 367315
rect 580981 365564 581227 366286
rect 583575 361027 584320 361051
rect 583575 360769 583603 361027
rect 584293 360769 584320 361027
rect 583575 360746 584320 360769
rect 290311 30949 290511 32541
rect 290073 30905 290992 30949
rect 290073 30361 290122 30905
rect 290933 30361 290992 30905
rect 290073 30317 290992 30361
<< via1 >>
rect 513911 593259 520276 609778
rect 556508 593934 560007 601770
rect 510907 570179 518330 576926
rect 556611 563187 560065 572886
rect 25460 486521 26354 500270
rect 20480 479565 20783 480450
rect 22005 480350 22308 481235
rect 21268 476599 21751 476743
rect 4728 470506 6108 475393
rect 19136 470495 24029 475286
rect 7486 467721 7690 468312
rect 7523 461352 8290 461984
rect 6476 438897 6728 439485
rect 7391 438204 7570 439002
rect 1738 435716 2398 435904
rect 13238 437442 14564 437642
rect 6378 429877 7086 430832
rect 4522 425868 4717 426541
rect 580981 366286 581227 367266
rect 583603 360769 584293 361027
rect 290122 30361 290933 30905
<< metal2 >>
rect 279035 644086 282907 644146
rect 279035 643726 282767 643786
rect 279035 554086 282627 554146
rect 279035 553726 282487 553786
rect 25311 500270 26552 500469
rect 25311 492593 25460 500270
rect 25262 486521 25460 492593
rect 26354 492593 26552 500270
rect 26354 492430 38581 492593
rect 26354 486659 28395 492430
rect 38334 486659 38581 492430
rect 26354 486521 38581 486659
rect 25262 486422 38581 486521
rect 25311 486372 26552 486422
rect 4420 475393 12415 475493
rect 4420 470506 4728 475393
rect 6108 470506 6256 475393
rect 4420 470365 6256 470506
rect 12269 470365 12415 475393
rect 4420 470219 12415 470365
rect 15695 469792 15851 482422
rect 15621 469755 15920 469792
rect 2247 469256 2511 469276
rect 2247 468578 2262 469256
rect 2494 468578 2511 469256
rect 7459 469236 8334 469270
rect 7459 469100 7494 469236
rect 8300 469100 8334 469236
rect 7459 469073 8334 469100
rect 15621 469083 15660 469755
rect 15889 469083 15920 469755
rect 2247 468557 2511 468578
rect 2268 461435 2475 468557
rect 7505 468354 7690 469073
rect 15621 469053 15920 469083
rect 7456 468312 7723 468354
rect 7456 467721 7486 468312
rect 7690 467721 7723 468312
rect 7456 467681 7723 467721
rect 16967 467330 17123 482466
rect 18306 479594 18658 482471
rect 21973 481235 22340 481278
rect 20445 480450 20812 480490
rect 18196 479537 18710 479594
rect 18196 478121 18241 479537
rect 18645 478121 18710 479537
rect 20445 479565 20480 480450
rect 20783 479975 20812 480450
rect 21973 480350 22005 481235
rect 22308 480747 22340 481235
rect 136829 481050 140840 481122
rect 136829 480747 136929 481050
rect 22308 480414 136929 480747
rect 140755 480747 140840 481050
rect 140755 480414 140936 480747
rect 22308 480350 140936 480414
rect 21973 480346 140936 480350
rect 21973 480310 22340 480346
rect 128830 479975 132831 479982
rect 20783 479922 140936 479975
rect 20783 479574 128886 479922
rect 20783 479565 20812 479574
rect 20445 479522 20812 479565
rect 128830 479271 128886 479574
rect 132750 479574 140936 479922
rect 132750 479271 132831 479574
rect 128830 479211 132831 479271
rect 18196 478064 18710 478121
rect 21251 476743 21774 476758
rect 21251 476599 21268 476743
rect 21751 476733 21774 476743
rect 21751 476633 142568 476733
rect 21751 476599 21774 476633
rect 21251 476583 21774 476599
rect 18828 475286 24285 475543
rect 18828 470495 19136 475286
rect 24029 470495 24285 475286
rect 18828 470214 24285 470495
rect 4524 467174 17123 467330
rect 1703 435904 2427 435927
rect 1703 435716 1738 435904
rect 2398 435889 2427 435904
rect 4524 435889 4680 467174
rect 7466 461984 8347 462028
rect 7466 461352 7523 461984
rect 8290 461352 8347 461984
rect 7466 461302 8347 461352
rect 5382 456631 5786 456990
rect 5343 456528 6129 456631
rect 5343 455115 5436 456528
rect 6072 455115 6129 456528
rect 10238 456434 10524 458058
rect 10720 457049 10842 458191
rect 10962 458053 140941 458106
rect 10962 457796 136913 458053
rect 136832 457377 136913 457796
rect 140759 457796 140941 458053
rect 140759 457377 140827 457796
rect 127385 457211 134893 457333
rect 136832 457317 140827 457377
rect 127385 457049 127507 457211
rect 10720 456927 127507 457049
rect 134771 456973 134893 457211
rect 128832 456791 132834 456858
rect 134771 456851 142279 456973
rect 128832 456434 128913 456791
rect 10238 456233 128913 456434
rect 132752 456233 132834 456791
rect 10238 456148 132834 456233
rect 5343 455031 6129 455115
rect 6463 439503 6744 439504
rect 6462 439485 6744 439503
rect 6462 438897 6476 439485
rect 6728 438897 6744 439485
rect 6462 438880 6744 438897
rect 6463 437005 6744 438880
rect 7368 439002 7592 439029
rect 7368 438204 7391 439002
rect 7570 438204 7592 439002
rect 7368 438178 7592 438204
rect 6447 436988 6755 437005
rect 6447 436151 6459 436988
rect 6743 436151 6755 436988
rect 6447 436136 6755 436151
rect 2398 435733 4680 435889
rect 2398 435716 2427 435733
rect 1703 435690 2427 435716
rect 7418 434511 7549 438178
rect 13208 437642 14598 437666
rect 13208 437442 13238 437642
rect 14564 437442 14598 437642
rect 13208 437416 14598 437442
rect 13394 436761 14363 437416
rect 13382 436724 14416 436761
rect 13382 434895 13424 436724
rect 14366 434895 14416 436724
rect 13382 434848 14416 434895
rect 7418 434380 141773 434511
rect 136831 434133 140827 434200
rect 136831 433676 136929 434133
rect 10249 433457 136929 433676
rect 140750 433676 140827 434133
rect 140750 433457 140833 433676
rect 10249 433366 140833 433457
rect 10219 433124 141383 433246
rect 10226 432924 132846 432928
rect 10226 432842 132847 432924
rect 10226 432642 128909 432842
rect 128832 432251 128909 432642
rect 132750 432251 132847 432842
rect 128832 432179 132847 432251
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 6302 429814 7162 429877
rect 11637 428240 13660 428297
rect 11637 428190 11697 428240
rect 11379 427828 11697 428190
rect 13585 428190 13660 428240
rect 13585 427828 13661 428190
rect 11379 427786 13661 427828
rect 11637 427782 13660 427786
rect 4524 426575 4680 426577
rect 4484 426541 4759 426575
rect 4484 425868 4522 426541
rect 4717 425868 4759 426541
rect 4484 425830 4759 425868
rect 3425 360329 135815 360419
rect 3425 350850 3515 360329
rect 3711 359987 135473 360077
rect 3711 351650 3801 359987
rect 4063 359639 135125 359729
rect 4063 352450 4153 359639
rect 52370 359282 134778 359382
rect 52370 357580 52470 359282
rect 51740 357480 52470 357580
rect 52658 358928 134424 359028
rect 52658 356580 52758 358928
rect 51612 356480 52758 356580
rect 53062 358592 134088 358692
rect 53062 355580 53162 358592
rect 51612 355480 53162 355580
rect 53382 358220 133716 358320
rect 53382 354580 53482 358220
rect 51636 354480 53482 354580
rect 53680 357796 133292 357896
rect 53680 353580 53780 357796
rect 51702 353480 53780 353580
rect 53946 357476 132972 357576
rect 53946 352580 54046 357476
rect 51736 352480 54046 352580
rect 4063 352360 5233 352450
rect 3711 351560 5211 351650
rect 3425 350760 5111 350850
rect 72760 283860 73112 283872
rect 72760 283841 72774 283860
rect 69998 283777 72774 283841
rect 72760 283754 72774 283777
rect 73100 283754 73112 283860
rect 72760 283742 73112 283754
rect 74040 279771 74668 279784
rect 74040 279756 74063 279771
rect 69640 279692 74063 279756
rect 74040 279659 74063 279692
rect 74651 279659 74668 279771
rect 74040 279641 74668 279659
rect 69609 267871 74311 267937
rect 69615 267216 74320 267280
rect 69642 265310 74369 265370
rect 70000 264731 132372 264791
rect 69965 264231 131889 264291
rect 69637 263773 131631 263833
rect 126401 249346 126485 249530
rect 126317 249334 126591 249346
rect 126317 249227 126333 249334
rect 126572 249227 126591 249334
rect 126317 249215 126591 249227
rect 66970 148120 67388 148132
rect 66970 148095 66984 148120
rect 62972 148043 66984 148095
rect 66970 148022 66984 148043
rect 67376 148022 67388 148120
rect 66970 148010 67388 148022
rect 66865 143880 67308 143889
rect 66865 143872 66876 143880
rect 62988 143808 66876 143872
rect 66865 143790 66876 143808
rect 67297 143790 67308 143880
rect 66865 143780 67308 143790
rect 46234 113554 124905 113564
rect 46234 113496 46264 113554
rect 46461 113496 124905 113554
rect 46234 113489 124905 113496
rect 46234 113356 124705 113364
rect 46234 113298 47992 113356
rect 48189 113298 124705 113356
rect 46234 113289 124705 113298
rect 46234 113154 124505 113164
rect 46234 113096 49795 113154
rect 49992 113096 124505 113154
rect 46234 113089 124505 113096
rect 46234 112956 124305 112964
rect 46234 112898 50047 112956
rect 50244 112898 124305 112956
rect 46234 112889 124305 112898
rect 46234 112755 124105 112764
rect 46234 112697 50335 112755
rect 50532 112697 124105 112755
rect 46234 112689 124105 112697
rect 46234 112554 123905 112564
rect 46234 112496 50615 112554
rect 50812 112496 123905 112554
rect 46234 112489 123905 112496
rect 79021 78218 79536 78232
rect 79021 78187 79036 78218
rect 74898 78123 79036 78187
rect 79021 78016 79036 78123
rect 79518 78016 79536 78218
rect 79021 77998 79536 78016
rect 79030 74215 79584 74230
rect 74562 74187 74618 74196
rect 79030 74187 79047 74215
rect 74545 74123 74554 74187
rect 74618 74123 79047 74187
rect 74562 74114 74618 74123
rect 79030 74075 79047 74123
rect 79566 74075 79584 74215
rect 79030 74060 79584 74075
rect 74987 56758 76924 56786
rect 74994 56114 76329 56142
rect 74982 50318 76028 50346
rect 76000 45421 76028 50318
rect 76300 45609 76328 56114
rect 76896 45818 76924 56758
rect 76896 45790 123222 45818
rect 76300 45581 123000 45609
rect 76000 45393 122769 45421
rect 56809 45168 122556 45175
rect 56809 45109 56820 45168
rect 57027 45109 122556 45168
rect 56809 45099 122556 45109
rect 56809 44966 122356 44975
rect 56809 44907 57406 44966
rect 57613 44907 122356 44966
rect 56809 44899 122356 44907
rect 56809 44767 122156 44775
rect 56809 44708 59488 44767
rect 59695 44708 122156 44767
rect 56809 44699 122156 44708
rect 56809 44567 121956 44575
rect 56809 44508 59793 44567
rect 60000 44508 121956 44567
rect 56809 44499 121956 44508
rect 56809 44367 121756 44375
rect 56809 44308 60146 44367
rect 60353 44308 121756 44367
rect 56809 44299 121756 44308
rect 56809 44167 121556 44175
rect 56809 44108 63928 44167
rect 64135 44108 121556 44167
rect 56809 44099 121556 44108
rect 56809 43967 121356 43975
rect 56809 43908 65290 43967
rect 65497 43908 121356 43967
rect 56809 43899 121356 43908
rect 56809 43767 121156 43775
rect 56809 43708 67318 43767
rect 67525 43708 121156 43767
rect 56809 43699 121156 43708
rect 121080 10348 121156 43699
rect 121107 4783 121156 10348
rect 121280 4983 121356 43899
rect 121480 5183 121556 44099
rect 121680 5383 121756 44299
rect 121880 5583 121956 44499
rect 122080 5783 122156 44699
rect 122280 5983 122356 44899
rect 122480 6183 122556 45099
rect 122741 6468 122769 45393
rect 122972 6725 123000 45581
rect 123194 6947 123222 45790
rect 123830 7371 123905 112489
rect 124030 7571 124105 112689
rect 124230 7771 124305 112889
rect 124430 7971 124505 113089
rect 124630 8171 124705 113289
rect 124830 8371 124905 113489
rect 126401 8765 126485 249215
rect 126801 249083 126885 249530
rect 126734 249073 127008 249083
rect 126734 248966 126750 249073
rect 126989 248966 127008 249073
rect 126734 248952 127008 248966
rect 126801 9110 126885 248952
rect 127201 248782 127285 249530
rect 127121 248773 127395 248782
rect 127121 248666 127136 248773
rect 127375 248666 127395 248773
rect 127121 248651 127395 248666
rect 127201 9455 127285 248651
rect 127601 248460 127685 249530
rect 127538 248447 127812 248460
rect 127538 248340 127557 248447
rect 127796 248340 127812 248447
rect 127538 248329 127812 248340
rect 127601 9786 127685 248329
rect 128001 248162 128085 249530
rect 127915 248150 128189 248162
rect 127915 248043 127934 248150
rect 128173 248043 128189 248150
rect 127915 248031 128189 248043
rect 128001 10175 128085 248031
rect 131571 10413 131631 263773
rect 131829 10717 131889 264231
rect 132312 11042 132372 264731
rect 132872 11398 132972 357476
rect 133192 11794 133292 357796
rect 133616 12132 133716 358220
rect 133988 12472 134088 358592
rect 134324 12866 134424 358928
rect 134678 13348 134778 359282
rect 135035 13783 135125 359639
rect 135383 14233 135473 359987
rect 135725 14607 135815 360329
rect 141261 15423 141383 433124
rect 141642 15813 141773 434380
rect 142157 16319 142279 456851
rect 142468 16608 142568 476633
rect 279035 464086 282347 464146
rect 279035 463726 282207 463786
rect 279035 374086 282067 374146
rect 279035 373726 281927 373786
rect 279035 284086 281787 284146
rect 279035 283726 281647 283786
rect 279035 194086 281507 194146
rect 279035 193726 281367 193786
rect 279035 104086 281227 104146
rect 279035 103726 281087 103786
rect 142468 16508 259100 16608
rect 142157 16197 255583 16319
rect 141642 15682 252014 15813
rect 141261 15301 248471 15423
rect 135725 14517 244917 14607
rect 135383 14143 241381 14233
rect 135035 13693 237833 13783
rect 134678 13248 234278 13348
rect 134324 12766 230730 12866
rect 133988 12372 227204 12472
rect 133616 12032 223656 12132
rect 133192 11694 220118 11794
rect 132872 11298 216560 11398
rect 132312 10982 212993 11042
rect 131829 10657 209466 10717
rect 131571 10353 205925 10413
rect 128001 10091 202384 10175
rect 128001 10085 128085 10091
rect 127601 9702 198829 9786
rect 127201 9371 195265 9455
rect 126801 9026 191710 9110
rect 126401 8681 188165 8765
rect 124830 8296 184626 8371
rect 124630 8096 181071 8171
rect 124430 7896 177531 7971
rect 124230 7696 173990 7771
rect 124030 7496 170464 7571
rect 123830 7296 166895 7371
rect 123194 6919 163320 6947
rect 122972 6697 159770 6725
rect 122741 6440 156252 6468
rect 122480 6107 152703 6183
rect 122280 5907 149162 5983
rect 122080 5707 145621 5783
rect 121880 5507 142052 5583
rect 121680 5307 138540 5383
rect 121480 5107 134985 5183
rect 121280 4907 131430 4983
rect 121107 4734 127890 4783
rect 127841 1280 127890 4734
rect 131354 1280 131430 4907
rect 134909 1280 134985 5107
rect 138464 1280 138540 5307
rect 141976 1280 142052 5507
rect 145545 1280 145621 5707
rect 149086 1280 149162 5907
rect 152627 1280 152703 6107
rect 156224 1280 156252 6440
rect 159742 1280 159770 6697
rect 163292 1280 163320 6919
rect 1324 800 1436 1280
rect 2506 800 2618 1280
rect 3688 800 3800 1280
rect 4870 800 4982 1280
rect 6052 800 6164 1280
rect 7234 800 7346 1280
rect 8416 800 8528 1280
rect 9598 800 9710 1280
rect 10780 800 10892 1280
rect 11962 800 12074 1280
rect 13144 800 13256 1280
rect 14326 800 14438 1280
rect 15508 800 15620 1280
rect 16690 800 16802 1280
rect 17872 800 17984 1280
rect 19054 800 19166 1280
rect 20236 800 20348 1280
rect 21418 800 21530 1280
rect 22600 800 22712 1280
rect 23782 800 23894 1280
rect 24964 800 25076 1280
rect 26146 800 26258 1280
rect 27328 800 27440 1280
rect 28510 800 28622 1280
rect 29692 800 29804 1280
rect 30874 800 30986 1280
rect 32056 800 32168 1280
rect 33238 800 33350 1280
rect 34420 800 34532 1280
rect 35602 800 35714 1280
rect 36784 800 36896 1280
rect 37966 800 38078 1280
rect 39148 800 39260 1280
rect 40330 800 40442 1280
rect 41512 800 41624 1280
rect 42694 800 42806 1280
rect 43876 800 43988 1280
rect 45058 800 45170 1280
rect 46240 800 46352 1280
rect 47422 800 47534 1280
rect 48604 800 48716 1280
rect 49786 800 49898 1280
rect 50968 800 51080 1280
rect 52150 800 52262 1280
rect 53332 800 53444 1280
rect 54514 800 54626 1280
rect 55696 800 55808 1280
rect 56878 800 56990 1280
rect 58060 800 58172 1280
rect 59242 800 59354 1280
rect 60424 800 60536 1280
rect 61606 800 61718 1280
rect 62788 800 62900 1280
rect 63970 800 64082 1280
rect 65152 800 65264 1280
rect 66334 800 66446 1280
rect 67516 800 67628 1280
rect 68698 800 68810 1280
rect 69880 800 69992 1280
rect 71062 800 71174 1280
rect 72244 800 72356 1280
rect 73426 800 73538 1280
rect 74608 800 74720 1280
rect 75790 800 75902 1280
rect 76972 800 77084 1280
rect 78154 800 78266 1280
rect 79336 800 79448 1280
rect 80518 800 80630 1280
rect 81700 800 81812 1280
rect 82882 800 82994 1280
rect 84064 800 84176 1280
rect 85246 800 85358 1280
rect 86428 800 86540 1280
rect 87610 800 87722 1280
rect 88792 800 88904 1280
rect 89974 800 90086 1280
rect 91156 800 91268 1280
rect 92338 800 92450 1280
rect 93520 800 93632 1280
rect 94702 800 94814 1280
rect 95884 800 95996 1280
rect 97066 800 97178 1280
rect 98248 800 98360 1280
rect 99430 800 99542 1280
rect 100612 800 100724 1280
rect 101794 800 101906 1280
rect 102976 800 103088 1280
rect 104158 800 104270 1280
rect 105340 800 105452 1280
rect 106522 800 106634 1280
rect 107704 800 107816 1280
rect 108886 800 108998 1280
rect 110068 800 110180 1279
rect 111250 800 111362 1280
rect 112432 800 112544 1280
rect 113614 800 113726 1280
rect 114796 800 114908 1280
rect 115978 800 116090 1280
rect 117160 800 117272 1280
rect 118342 800 118454 1280
rect 119524 800 119636 1280
rect 120706 800 120818 1280
rect 121888 800 122000 1280
rect 123070 800 123182 1280
rect 124252 800 124364 1280
rect 125434 800 125546 1280
rect 126616 800 126728 1280
rect 127798 800 127910 1280
rect 128980 800 129092 1280
rect 130162 800 130274 1280
rect 131344 800 131456 1280
rect 132526 800 132638 1280
rect 133708 800 133820 1280
rect 134890 800 135002 1280
rect 136072 800 136184 1280
rect 137254 800 137366 1280
rect 138479 1279 138528 1280
rect 141992 1279 142068 1280
rect 145547 1279 145623 1280
rect 149102 1279 149178 1280
rect 152614 1279 152690 1280
rect 156183 1279 156259 1280
rect 159724 1279 159800 1280
rect 163265 1279 163341 1280
rect 166820 1279 166895 7296
rect 170389 1279 170464 7496
rect 173915 1279 173990 7696
rect 177456 1279 177531 7896
rect 180996 1279 181071 8096
rect 184551 1279 184626 8296
rect 188081 1280 188165 8681
rect 191626 1280 191710 9026
rect 195181 8597 195265 9371
rect 198745 8942 198829 9702
rect 202300 9287 202384 10091
rect 195181 1280 195268 8597
rect 198736 1280 198829 8942
rect 202287 9138 202384 9287
rect 205846 9812 205925 10353
rect 202287 1280 202371 9138
rect 205846 1280 205930 9812
rect 209382 1280 209466 10657
rect 212933 1280 212993 10982
rect 216460 1280 216560 11298
rect 220018 1280 220118 11694
rect 223556 1280 223656 12032
rect 227104 1280 227204 12372
rect 230630 1280 230730 12766
rect 234178 1280 234278 13248
rect 237743 1280 237833 13693
rect 241291 1280 241381 14143
rect 244827 1280 244917 14517
rect 248349 1280 248471 15301
rect 251883 1280 252014 15682
rect 255461 1280 255583 16197
rect 259000 1280 259100 16508
rect 262274 9685 262334 11294
rect 265822 9812 265882 11294
rect 269370 9942 269430 11294
rect 272918 10070 272978 11294
rect 276466 10196 276526 11294
rect 278214 10324 278274 11294
rect 278562 10452 278622 11294
rect 278910 10582 278970 11294
rect 279258 10709 279318 11294
rect 279606 10837 279666 11294
rect 279954 10965 280014 11294
rect 280302 11093 280362 11294
rect 280227 11088 280448 11093
rect 280227 11032 280236 11088
rect 280439 11032 280448 11088
rect 280227 11027 280448 11032
rect 279879 10960 280100 10965
rect 279879 10904 279888 10960
rect 280091 10904 280100 10960
rect 279879 10899 280100 10904
rect 279510 10832 279731 10837
rect 279510 10776 279573 10832
rect 279722 10776 279731 10832
rect 279510 10771 279731 10776
rect 279186 10704 279407 10709
rect 279186 10648 279262 10704
rect 279398 10648 279407 10704
rect 279186 10643 279407 10648
rect 278837 10577 279058 10582
rect 278837 10521 278859 10577
rect 279049 10521 279058 10577
rect 278837 10516 279058 10521
rect 278479 10447 278700 10452
rect 278479 10391 278570 10447
rect 278691 10391 278700 10447
rect 278479 10386 278700 10391
rect 278145 10319 278366 10324
rect 278145 10263 278154 10319
rect 278357 10263 278366 10319
rect 278145 10258 278366 10263
rect 276390 10191 276611 10196
rect 276390 10135 276399 10191
rect 276602 10135 276611 10191
rect 276390 10130 276611 10135
rect 272836 10065 273050 10070
rect 272836 10009 272845 10065
rect 273048 10009 273050 10065
rect 272836 10004 273050 10009
rect 269312 9937 269533 9942
rect 269312 9881 269321 9937
rect 269524 9881 269533 9937
rect 269312 9876 269533 9881
rect 265735 9807 265956 9812
rect 265735 9751 265744 9807
rect 265947 9751 265956 9807
rect 265735 9746 265956 9751
rect 262190 9680 262411 9685
rect 262190 9624 262199 9680
rect 262402 9624 262411 9680
rect 262190 9619 262411 9624
rect 262274 7841 262334 9619
rect 265822 8091 265882 9746
rect 269370 8330 269430 9876
rect 272918 8569 272978 10004
rect 276466 8842 276526 10130
rect 276466 8782 276809 8842
rect 272918 8509 273261 8569
rect 269370 8270 269714 8330
rect 265822 8031 266178 8091
rect 262274 7781 262630 7841
rect 262570 1280 262630 7781
rect 266118 1280 266178 8031
rect 269654 1280 269714 8270
rect 273201 1280 273261 8509
rect 276749 1280 276809 8782
rect 278214 3103 278274 10258
rect 278562 3410 278622 10386
rect 278910 3660 278970 10516
rect 279258 3967 279318 10643
rect 279606 4320 279666 10771
rect 279954 4581 280014 10899
rect 280302 4820 280362 11027
rect 281027 5033 281087 103726
rect 281167 5173 281227 104086
rect 281307 5313 281367 193726
rect 281447 5453 281507 194086
rect 281587 5593 281647 283726
rect 281727 5733 281787 284086
rect 281867 5873 281927 373726
rect 282007 6013 282067 374086
rect 282147 6153 282207 463726
rect 282287 6293 282347 464086
rect 282427 6433 282487 553726
rect 282567 6573 282627 554086
rect 282707 6713 282767 643726
rect 282847 6853 282907 644086
rect 303822 644086 307687 644146
rect 286531 277791 286590 277827
rect 286531 9685 286590 277613
rect 298623 277776 298693 277829
rect 286731 277121 286790 277195
rect 286731 9813 286790 276926
rect 286931 275993 286990 276086
rect 286931 9941 286990 275798
rect 287131 273905 287190 273992
rect 287131 10069 287190 273710
rect 287331 271810 287390 271952
rect 287331 10198 287390 271615
rect 287531 269719 287590 269792
rect 287531 10325 287590 269524
rect 287731 266547 287790 266628
rect 287731 10453 287790 266352
rect 287931 261294 287990 261356
rect 287931 10581 287990 261087
rect 298423 260788 298493 260847
rect 298223 208190 298293 208297
rect 288131 197629 288190 197695
rect 288131 10709 288190 197431
rect 298023 155592 298093 155657
rect 297823 102990 297893 103167
rect 288309 87181 288390 87208
rect 288309 86937 288390 86979
rect 288331 10837 288390 86937
rect 288552 79455 288870 79519
rect 288552 10965 288616 79455
rect 297472 47527 297693 47597
rect 288910 47431 289456 47493
rect 288910 11093 288972 47431
rect 297246 46310 297494 46449
rect 290073 30905 290992 30949
rect 290073 30361 290122 30905
rect 290933 30361 290992 30905
rect 290073 30317 290992 30361
rect 288826 11088 289047 11093
rect 288826 11032 288835 11088
rect 289038 11032 289047 11088
rect 288826 11027 289047 11032
rect 288452 10960 288673 10965
rect 288452 10904 288461 10960
rect 288664 10904 288673 10960
rect 288452 10899 288673 10904
rect 288248 10832 288469 10837
rect 288248 10776 288257 10832
rect 288460 10776 288469 10832
rect 288248 10771 288469 10776
rect 288053 10704 288274 10709
rect 288053 10648 288062 10704
rect 288265 10648 288274 10704
rect 288053 10643 288274 10648
rect 287856 10576 288077 10581
rect 287856 10520 287865 10576
rect 288068 10520 288077 10576
rect 287856 10515 288077 10520
rect 287654 10448 287875 10453
rect 287654 10392 287663 10448
rect 287866 10392 287875 10448
rect 287654 10387 287875 10392
rect 287455 10320 287676 10325
rect 287455 10264 287464 10320
rect 287667 10264 287676 10320
rect 287455 10259 287676 10264
rect 287246 10193 287467 10198
rect 287246 10137 287255 10193
rect 287458 10137 287467 10193
rect 287246 10132 287467 10137
rect 287060 10064 287281 10069
rect 287060 10008 287069 10064
rect 287272 10008 287281 10064
rect 287060 10003 287281 10008
rect 286857 9936 287078 9941
rect 286857 9880 286866 9936
rect 287069 9880 287078 9936
rect 286857 9875 287078 9880
rect 286670 9808 286891 9813
rect 286670 9752 286679 9808
rect 286882 9752 286891 9808
rect 286670 9747 286891 9752
rect 286452 9680 286673 9685
rect 286452 9624 286461 9680
rect 286664 9624 286673 9680
rect 286452 9619 286673 9624
rect 286531 9520 286590 9619
rect 286731 9520 286790 9747
rect 286931 9520 286990 9875
rect 287131 9520 287190 10003
rect 287331 9520 287390 10132
rect 287531 9520 287590 10259
rect 287731 9520 287790 10387
rect 287931 9520 287990 10515
rect 288131 9520 288190 10643
rect 288331 9520 288390 10771
rect 288552 9520 288616 10899
rect 288910 9520 288972 11027
rect 297423 10535 297493 46310
rect 297350 10530 297571 10535
rect 297350 10474 297359 10530
rect 297562 10474 297571 10530
rect 297350 10469 297571 10474
rect 297423 9617 297493 10469
rect 297623 10407 297693 47527
rect 297546 10402 297767 10407
rect 297546 10346 297555 10402
rect 297758 10346 297767 10402
rect 297546 10341 297767 10346
rect 297623 9617 297693 10341
rect 297823 10279 297893 102785
rect 297744 10274 297965 10279
rect 297744 10218 297753 10274
rect 297956 10218 297965 10274
rect 297744 10213 297965 10218
rect 297823 9617 297893 10213
rect 298023 10150 298093 155388
rect 297951 10145 298172 10150
rect 297951 10089 297960 10145
rect 298163 10089 298172 10145
rect 297951 10084 298172 10089
rect 298023 9617 298093 10084
rect 298223 10023 298293 207988
rect 298149 10018 298370 10023
rect 298149 9962 298158 10018
rect 298361 9962 298370 10018
rect 298149 9957 298370 9962
rect 298223 9617 298293 9957
rect 298423 9895 298493 260587
rect 298345 9890 298566 9895
rect 298345 9834 298354 9890
rect 298557 9834 298566 9890
rect 298345 9829 298566 9834
rect 298423 9617 298493 9829
rect 298623 9767 298693 277538
rect 298541 9762 298762 9767
rect 298541 9706 298550 9762
rect 298753 9706 298762 9762
rect 298541 9701 298762 9706
rect 298623 9617 298693 9701
rect 303822 7132 303882 644086
rect 303962 643726 307687 643786
rect 303962 7352 304022 643726
rect 444175 617823 448174 617824
rect 444175 617699 560181 617823
rect 444175 614087 444372 617699
rect 448011 614087 560181 617699
rect 444175 613931 560181 614087
rect 444223 613929 560181 613931
rect 513415 609778 520733 610315
rect 513415 593259 513911 609778
rect 520276 593259 520733 609778
rect 556287 602040 560181 613929
rect 556287 601770 560183 602040
rect 556287 593934 556508 601770
rect 560007 593934 560183 601770
rect 556287 593698 560183 593934
rect 513415 592789 520733 593259
rect 583563 589372 583751 589414
rect 583563 588859 583568 589372
rect 583746 588859 583751 589372
rect 583563 588791 583751 588859
rect 583568 587366 583746 588791
rect 563565 587188 583746 587366
rect 563548 582534 565009 582654
rect 510422 576926 518844 577547
rect 510422 570179 510907 576926
rect 518330 570179 518844 576926
rect 510422 569612 518844 570179
rect 556374 572886 560268 573078
rect 556374 566873 556611 572886
rect 452076 566724 556611 566873
rect 452076 563112 452351 566724
rect 455990 563187 556611 566724
rect 560065 566873 560268 572886
rect 560065 563187 560278 566873
rect 455990 563112 560278 563187
rect 452076 562979 560278 563112
rect 438929 561647 439466 561660
rect 438929 561526 438947 561647
rect 439446 561643 439466 561647
rect 564895 561643 565009 582534
rect 439446 561529 565009 561643
rect 439446 561526 439466 561529
rect 438929 561509 439466 561526
rect 304102 554086 307687 554146
rect 304102 7561 304162 554086
rect 304242 553726 307687 553786
rect 304242 7746 304302 553726
rect 304382 464086 307687 464146
rect 304382 7899 304442 464086
rect 304522 463726 307687 463786
rect 304522 8078 304582 463726
rect 557755 435818 557986 435844
rect 557755 434769 557782 435818
rect 557961 434975 557986 435818
rect 557961 434769 559425 434975
rect 557755 434744 559425 434769
rect 582171 433815 583321 434170
rect 583433 433815 583444 434170
rect 582185 431416 583313 431771
rect 583425 431416 583453 431771
rect 423480 422228 425176 422253
rect 423480 422017 423509 422228
rect 425145 422188 425176 422228
rect 425145 422035 559381 422188
rect 425145 422017 425176 422035
rect 423480 421993 425176 422017
rect 452250 421269 559235 421330
rect 452250 421117 452329 421269
rect 452172 420738 452329 421117
rect 452250 420650 452329 420738
rect 456074 421117 559235 421269
rect 456074 420738 559442 421117
rect 456074 420650 559235 420738
rect 452250 420572 559235 420650
rect 444312 419339 559230 419413
rect 444312 419211 444386 419339
rect 444073 418832 444386 419211
rect 444312 418708 444386 418832
rect 447969 419211 559230 419339
rect 447969 418832 559373 419211
rect 447969 418708 559230 418832
rect 444312 418647 559230 418708
rect 456842 415208 559384 415328
rect 304662 374086 307687 374146
rect 304662 8238 304722 374086
rect 304802 373726 307687 373786
rect 304802 8398 304862 373726
rect 304942 284086 307687 284146
rect 304942 8551 305002 284086
rect 305082 283726 307687 283786
rect 305082 8711 305142 283726
rect 305222 194086 307687 194146
rect 305222 8890 305282 194086
rect 305362 193726 307687 193786
rect 305362 9043 305422 193726
rect 305502 104086 307687 104146
rect 305502 9209 305562 104086
rect 305642 103726 307687 103786
rect 305642 9401 305702 103726
rect 404410 10535 404470 10715
rect 404329 10530 404550 10535
rect 404329 10474 404338 10530
rect 404541 10474 404550 10530
rect 404329 10469 404550 10474
rect 305642 9341 400929 9401
rect 305502 9149 397403 9209
rect 305362 8983 393845 9043
rect 305222 8830 390293 8890
rect 305082 8651 386748 8711
rect 304942 8491 383209 8551
rect 304802 8338 379657 8398
rect 304662 8178 376111 8238
rect 304522 8018 372540 8078
rect 304382 7839 369021 7899
rect 304242 7686 365456 7746
rect 304102 7501 361904 7561
rect 303962 7292 358382 7352
rect 303822 7072 354827 7132
rect 282847 6793 351281 6853
rect 282707 6653 347753 6713
rect 282567 6513 344193 6573
rect 282427 6373 340644 6433
rect 282287 6233 337105 6293
rect 282147 6093 333556 6153
rect 282007 5953 329996 6013
rect 281867 5813 326457 5873
rect 281727 5673 322918 5733
rect 281587 5533 319369 5593
rect 281447 5393 315830 5453
rect 281307 5253 312270 5313
rect 281167 5113 308742 5173
rect 281027 4973 305182 5033
rect 280302 4760 301629 4820
rect 279954 4521 298093 4581
rect 279606 4260 294546 4320
rect 279258 3907 290998 3967
rect 278910 3600 287451 3660
rect 278562 3350 283903 3410
rect 278214 3043 280356 3103
rect 280296 1280 280356 3043
rect 283843 1280 283903 3350
rect 287391 1280 287451 3600
rect 290938 1280 290998 3907
rect 294486 1280 294546 4260
rect 298033 1280 298093 4521
rect 301569 1280 301629 4760
rect 305122 1280 305182 4973
rect 308682 1280 308742 5113
rect 312210 1280 312270 5253
rect 315770 1280 315830 5393
rect 319309 1280 319369 5533
rect 322858 1280 322918 5673
rect 326397 1280 326457 5813
rect 329936 1280 329996 5953
rect 333496 1280 333556 6093
rect 337045 1280 337105 6233
rect 340584 1280 340644 6373
rect 344133 1280 344193 6513
rect 347693 1280 347753 6653
rect 351221 1280 351281 6793
rect 354767 1280 354827 7072
rect 358322 1280 358382 7292
rect 361844 1280 361904 7501
rect 365396 1634 365456 7686
rect 368961 1280 369021 7839
rect 372480 1280 372540 8018
rect 376051 1280 376111 8178
rect 379597 1280 379657 8338
rect 383149 1280 383209 8491
rect 386688 1280 386748 8651
rect 390233 1280 390293 8830
rect 393785 1280 393845 8983
rect 397343 1280 397403 9149
rect 400869 1280 400929 9341
rect 404410 1280 404470 10469
rect 407958 10407 408018 10715
rect 407883 10402 408104 10407
rect 407883 10346 407892 10402
rect 408095 10346 408104 10402
rect 407883 10341 408104 10346
rect 407958 1280 408018 10341
rect 411506 10279 411566 10715
rect 411441 10274 411662 10279
rect 411441 10218 411450 10274
rect 411653 10218 411662 10274
rect 411441 10213 411662 10218
rect 411506 1280 411566 10213
rect 415054 10149 415114 10667
rect 414989 10144 415210 10149
rect 414989 10088 414998 10144
rect 415201 10088 415210 10144
rect 414989 10083 415210 10088
rect 415054 1280 415114 10083
rect 418602 10022 418662 10667
rect 418526 10017 418747 10022
rect 418526 9961 418535 10017
rect 418738 9961 418747 10017
rect 418526 9956 418747 9961
rect 418602 1280 418662 9956
rect 422150 9893 422210 10667
rect 422062 9888 422283 9893
rect 422062 9832 422071 9888
rect 422274 9832 422283 9888
rect 422062 9827 422283 9832
rect 422150 1280 422210 9827
rect 425698 9766 425758 10667
rect 425636 9761 425857 9766
rect 425636 9705 425645 9761
rect 425848 9705 425857 9761
rect 425636 9700 425857 9705
rect 425698 1280 425758 9700
rect 456842 7086 456962 415208
rect 429205 6966 456962 7086
rect 457161 414489 559390 414609
rect 138436 800 138548 1279
rect 139618 800 139730 1279
rect 140800 800 140912 1279
rect 141982 800 142094 1279
rect 143164 800 143276 1279
rect 144346 800 144458 1279
rect 145528 1178 145648 1279
rect 145528 800 145640 1178
rect 146710 800 146822 1279
rect 147892 800 148004 1279
rect 149074 800 149186 1279
rect 150256 800 150368 1279
rect 151438 800 151550 1279
rect 152614 1096 152732 1279
rect 152620 800 152732 1096
rect 153802 800 153914 1279
rect 154984 800 155096 1279
rect 156166 800 156278 1279
rect 157348 800 157460 1279
rect 158530 800 158642 1279
rect 159712 1152 159836 1279
rect 159712 800 159824 1152
rect 160894 800 161006 1279
rect 162076 800 162188 1279
rect 163258 1108 163374 1279
rect 163258 800 163370 1108
rect 164440 800 164552 1279
rect 165622 800 165734 1279
rect 166804 1140 166922 1279
rect 166804 800 166916 1140
rect 167986 800 168098 1279
rect 169168 800 169280 1279
rect 170348 1130 170464 1279
rect 170350 1112 170464 1130
rect 170350 800 170462 1112
rect 171532 800 171644 1279
rect 172714 800 172826 1279
rect 173896 800 174008 1279
rect 175078 800 175190 1279
rect 176260 800 176372 1279
rect 177442 800 177554 1279
rect 178624 800 178736 1279
rect 179806 800 179918 1279
rect 180988 800 181100 1279
rect 182170 800 182282 1279
rect 183352 800 183464 1279
rect 184534 800 184646 1279
rect 185716 800 185828 1279
rect 186898 800 187010 1279
rect 188080 800 188192 1279
rect 189262 800 189374 1279
rect 190444 800 190556 1279
rect 191626 983 191738 1279
rect 191613 982 191738 983
rect 191626 800 191738 982
rect 192808 800 192920 1279
rect 193990 800 194102 1279
rect 195172 800 195284 1279
rect 196354 800 196466 1279
rect 197536 800 197648 1279
rect 198718 800 198830 1280
rect 199900 800 200012 1280
rect 201082 800 201194 1280
rect 202264 800 202376 1280
rect 203446 800 203558 1280
rect 204628 800 204740 1280
rect 205810 1279 205930 1280
rect 205810 800 205922 1279
rect 206992 800 207104 1280
rect 208174 800 208286 1280
rect 209356 800 209468 1280
rect 210538 800 210650 1280
rect 211720 800 211832 1280
rect 212902 800 213014 1280
rect 214084 800 214196 1280
rect 215266 800 215378 1280
rect 216448 800 216560 1280
rect 217630 800 217742 1280
rect 218812 800 218924 1280
rect 219994 1279 220118 1280
rect 219994 800 220106 1279
rect 221176 800 221288 1280
rect 222358 800 222470 1280
rect 223540 1279 223656 1280
rect 223540 800 223652 1279
rect 224722 800 224834 1280
rect 225904 800 226016 1280
rect 227086 1279 227204 1280
rect 227086 800 227198 1279
rect 228268 800 228380 1280
rect 229450 800 229562 1280
rect 230630 1279 230744 1280
rect 230632 800 230744 1279
rect 231814 800 231926 1280
rect 232996 800 233108 1280
rect 234178 800 234290 1280
rect 235360 800 235472 1280
rect 236542 800 236654 1280
rect 237724 800 237836 1280
rect 238906 800 239018 1280
rect 240088 800 240200 1280
rect 241270 800 241382 1280
rect 242452 800 242564 1280
rect 243634 800 243746 1280
rect 244816 800 244928 1280
rect 245998 800 246110 1280
rect 247180 800 247292 1280
rect 248362 800 248474 1280
rect 249544 800 249656 1280
rect 250726 800 250838 1280
rect 251908 800 252020 1280
rect 253090 800 253202 1280
rect 254272 800 254384 1280
rect 255454 800 255566 1280
rect 256636 800 256748 1280
rect 257818 800 257930 1280
rect 259000 800 259112 1280
rect 260182 800 260294 1280
rect 261364 800 261476 1280
rect 262546 800 262658 1280
rect 263728 800 263840 1280
rect 264910 800 265022 1280
rect 266092 800 266204 1280
rect 267274 800 267386 1280
rect 268456 800 268568 1280
rect 269638 1175 269752 1280
rect 269638 800 269750 1175
rect 270820 800 270932 1280
rect 272002 800 272114 1280
rect 273184 800 273296 1280
rect 274366 800 274478 1280
rect 275548 800 275660 1280
rect 276730 800 276842 1280
rect 277912 800 278024 1280
rect 279094 800 279206 1280
rect 280276 800 280388 1280
rect 281458 800 281570 1280
rect 282640 800 282752 1280
rect 283822 800 283934 1280
rect 285004 800 285116 1280
rect 286186 800 286298 1280
rect 287368 800 287480 1280
rect 288550 800 288662 1280
rect 289732 800 289844 1280
rect 290914 800 291026 1280
rect 292096 800 292208 1280
rect 293278 800 293390 1280
rect 294460 800 294572 1280
rect 295642 800 295754 1280
rect 296824 800 296936 1280
rect 298006 800 298118 1280
rect 299188 800 299300 1280
rect 300370 800 300482 1280
rect 301552 800 301664 1280
rect 302734 800 302846 1280
rect 303916 800 304028 1280
rect 305098 800 305210 1280
rect 306280 800 306392 1280
rect 307462 800 307574 1280
rect 308644 800 308756 1280
rect 309826 800 309938 1280
rect 311008 800 311120 1280
rect 312190 800 312302 1280
rect 313372 800 313484 1280
rect 314554 800 314666 1280
rect 315736 800 315848 1280
rect 316918 800 317030 1280
rect 318100 800 318212 1280
rect 319282 800 319394 1280
rect 320464 800 320576 1280
rect 321646 800 321758 1280
rect 322828 800 322940 1280
rect 324010 800 324122 1280
rect 325192 800 325304 1280
rect 326374 800 326486 1280
rect 327556 800 327668 1280
rect 328738 800 328850 1280
rect 329920 800 330032 1280
rect 331102 800 331214 1280
rect 332284 800 332396 1280
rect 333466 800 333578 1280
rect 334648 800 334760 1280
rect 335830 800 335942 1280
rect 337012 800 337124 1280
rect 338194 800 338306 1280
rect 339376 800 339488 1280
rect 340558 800 340670 1280
rect 341740 800 341852 1280
rect 342922 800 343034 1280
rect 344104 800 344216 1280
rect 345286 800 345398 1280
rect 346468 800 346580 1280
rect 347650 800 347762 1280
rect 348832 800 348944 1280
rect 350014 800 350126 1280
rect 351196 800 351308 1280
rect 352378 800 352490 1280
rect 353560 800 353672 1280
rect 354742 800 354854 1280
rect 355924 800 356036 1280
rect 357106 800 357218 1280
rect 358288 800 358400 1280
rect 359470 800 359582 1280
rect 360652 800 360764 1280
rect 361834 800 361946 1280
rect 363016 800 363128 1280
rect 364198 800 364310 1280
rect 365380 800 365492 1280
rect 366562 800 366674 1280
rect 367744 800 367856 1280
rect 368926 800 369038 1280
rect 370108 800 370220 1280
rect 371290 800 371402 1280
rect 372472 800 372584 1280
rect 373654 800 373766 1280
rect 374836 800 374948 1280
rect 376018 800 376130 1280
rect 377200 800 377312 1280
rect 378382 800 378494 1280
rect 379564 800 379676 1280
rect 380746 800 380858 1280
rect 381928 800 382040 1280
rect 383110 800 383222 1280
rect 384292 800 384404 1280
rect 385474 800 385586 1280
rect 386656 800 386768 1280
rect 387838 800 387950 1280
rect 389020 800 389132 1280
rect 390202 800 390314 1280
rect 391384 800 391496 1280
rect 392566 800 392678 1280
rect 393748 800 393860 1280
rect 394930 800 395042 1280
rect 396112 800 396224 1280
rect 397294 800 397406 1280
rect 398476 800 398588 1280
rect 399658 800 399770 1280
rect 400840 800 400952 1280
rect 402022 800 402134 1280
rect 403204 800 403316 1280
rect 404386 800 404498 1280
rect 405568 800 405680 1280
rect 406750 800 406862 1280
rect 407932 800 408044 1280
rect 409114 800 409226 1280
rect 410296 800 410408 1280
rect 411478 800 411590 1280
rect 412660 800 412772 1280
rect 413842 800 413954 1280
rect 415024 800 415136 1280
rect 416206 800 416318 1280
rect 417388 800 417500 1280
rect 418570 800 418682 1280
rect 419752 800 419864 1280
rect 420934 800 421046 1280
rect 422116 800 422228 1280
rect 423298 800 423410 1280
rect 424480 800 424592 1280
rect 425662 800 425774 1280
rect 426844 800 426956 1280
rect 428026 800 428138 1280
rect 429205 1176 429325 6966
rect 457161 6473 457281 414489
rect 547144 413369 559324 413371
rect 432738 6353 457281 6473
rect 458295 412900 458412 412928
rect 432738 1280 432858 6353
rect 458295 5617 458412 412283
rect 436289 5500 458412 5617
rect 458587 412900 458704 412934
rect 436289 1280 436406 5500
rect 458587 4993 458704 412283
rect 439839 4876 458704 4993
rect 458893 412900 459010 412937
rect 439839 1280 439956 4876
rect 458893 4549 459010 412283
rect 443388 4432 459010 4549
rect 459229 412900 459346 412930
rect 429208 800 429320 1176
rect 430390 800 430502 1280
rect 431572 800 431684 1280
rect 432738 1111 432866 1280
rect 432754 800 432866 1111
rect 433936 800 434048 1280
rect 435118 800 435230 1280
rect 436289 1014 436412 1280
rect 436300 800 436412 1014
rect 437482 800 437594 1280
rect 438664 800 438776 1280
rect 439839 981 439958 1280
rect 439846 800 439958 981
rect 441028 800 441140 1280
rect 442210 800 442322 1280
rect 443388 1014 443505 4432
rect 459229 3958 459346 412283
rect 446938 3841 459346 3958
rect 459597 412900 459714 412930
rect 547144 412928 547393 413369
rect 552551 412928 559324 413369
rect 466206 412763 473703 412769
rect 466196 412620 559318 412763
rect 466196 412320 466355 412620
rect 443392 800 443504 1014
rect 444574 800 444686 1280
rect 445756 800 445868 1280
rect 446938 1063 447055 3841
rect 459597 3448 459714 412283
rect 466206 410038 466355 412320
rect 473541 412320 559318 412620
rect 473541 410038 473703 412320
rect 466206 409865 473703 410038
rect 580930 369269 581274 369297
rect 580930 367739 580964 369269
rect 581233 367739 581274 369269
rect 580930 367703 581274 367739
rect 580981 367266 581227 367703
rect 580981 366233 581227 366286
rect 583575 361027 584320 361051
rect 583575 360769 583603 361027
rect 584293 360769 584320 361027
rect 583575 360746 584320 360769
rect 450488 3331 459714 3448
rect 450488 1280 450605 3331
rect 446938 800 447050 1063
rect 448120 800 448232 1280
rect 449302 800 449414 1280
rect 450484 1096 450605 1280
rect 450484 800 450596 1096
rect 451666 800 451778 1280
rect 452848 800 452960 1280
rect 454019 1122 454142 1280
rect 454030 800 454142 1122
rect 455212 800 455324 1280
rect 456394 800 456506 1280
rect 457576 1190 457696 1280
rect 457576 800 457688 1190
rect 458758 800 458870 1280
rect 459940 800 460052 1280
rect 461112 1086 461234 1280
rect 461122 800 461234 1086
rect 462304 800 462416 1280
rect 463486 800 463598 1280
rect 464668 1094 464787 1280
rect 464668 800 464780 1094
rect 465850 800 465962 1280
rect 467032 800 467144 1280
rect 468212 1163 468329 1280
rect 468214 800 468326 1163
rect 469396 800 469508 1280
rect 470578 800 470690 1280
rect 471754 1147 471872 1280
rect 471760 800 471872 1147
rect 472942 800 473054 1280
rect 474124 800 474236 1280
rect 475296 1117 475418 1280
rect 475306 800 475418 1117
rect 476488 800 476600 1280
rect 477670 800 477782 1280
rect 478852 800 478964 1280
rect 480034 800 480146 1280
rect 481216 800 481328 1280
rect 482398 800 482510 1280
rect 483580 800 483692 1280
rect 484762 800 484874 1280
rect 485944 800 486056 1280
rect 487126 800 487238 1280
rect 488308 800 488420 1280
rect 489490 800 489602 1280
rect 490672 800 490784 1280
rect 491854 800 491966 1280
rect 493036 800 493148 1280
rect 494218 800 494330 1280
rect 495400 800 495512 1280
rect 496582 800 496694 1280
rect 497764 800 497876 1280
rect 498946 800 499058 1280
rect 500128 800 500240 1280
rect 501310 800 501422 1280
rect 502492 800 502604 1280
rect 503674 800 503786 1280
rect 504856 800 504968 1280
rect 506038 800 506150 1280
rect 507220 800 507332 1280
rect 508402 800 508514 1280
rect 509584 800 509696 1280
rect 510766 800 510878 1280
rect 511948 800 512060 1280
rect 513130 800 513242 1280
rect 514312 800 514424 1280
rect 515494 800 515606 1280
rect 516676 800 516788 1280
rect 517858 800 517970 1280
rect 519040 800 519152 1280
rect 520222 800 520334 1280
rect 521404 800 521516 1280
rect 522586 800 522698 1280
rect 523768 800 523880 1280
rect 524950 800 525062 1280
rect 526132 800 526244 1280
rect 527314 800 527426 1280
rect 528496 800 528608 1280
rect 529678 800 529790 1280
rect 530860 800 530972 1280
rect 532042 800 532154 1280
rect 533224 800 533336 1280
rect 534406 800 534518 1280
rect 535588 800 535700 1280
rect 536770 800 536882 1280
rect 537952 800 538064 1280
rect 539134 800 539246 1280
rect 540316 800 540428 1280
rect 541498 800 541610 1280
rect 542680 800 542792 1280
rect 543862 800 543974 1280
rect 545044 800 545156 1280
rect 546226 800 546338 1280
rect 547408 800 547520 1280
rect 548590 800 548702 1280
rect 549772 800 549884 1280
rect 550954 800 551066 1280
rect 552136 800 552248 1280
rect 553318 800 553430 1280
rect 554500 800 554612 1280
rect 555682 800 555794 1280
rect 556864 800 556976 1280
rect 558046 800 558158 1280
rect 559228 800 559340 1280
rect 560410 800 560522 1280
rect 561592 800 561704 1280
rect 562774 800 562886 1280
rect 563956 800 564068 1280
rect 565138 800 565250 1280
rect 566320 800 566432 1280
rect 567502 800 567614 1280
rect 568684 800 568796 1280
rect 569866 800 569978 1280
rect 571048 800 571160 1280
rect 572230 800 572342 1280
rect 573412 800 573524 1280
rect 574594 800 574706 1280
rect 575776 800 575888 1280
rect 576958 800 577070 1280
rect 578140 800 578252 1280
rect 579322 800 579434 1280
rect 580504 800 580616 1280
rect 581686 800 581798 1280
rect 582868 800 582980 1280
rect 584050 800 584162 1280
rect 202266 0 202326 800
rect 205814 0 205874 800
rect 209362 0 209422 800
rect 212910 0 212970 800
rect 216458 0 216518 800
rect 220006 0 220066 800
rect 223554 0 223614 800
rect 227102 0 227162 800
rect 230650 0 230710 800
rect 234198 0 234258 800
rect 237746 0 237806 800
rect 241294 0 241354 800
rect 351222 0 351282 800
rect 354770 0 354830 800
rect 358318 0 358378 800
rect 361866 0 361926 800
rect 365414 0 365474 800
rect 368962 0 369022 800
<< via2 >>
rect 28395 486659 38334 492430
rect 6256 470365 12269 475393
rect 2262 468578 2494 469256
rect 7494 469100 8300 469236
rect 15660 469083 15889 469755
rect 18241 478121 18645 479537
rect 136929 480414 140755 481050
rect 128886 479271 132750 479922
rect 19136 470495 24029 475286
rect 7523 461352 8290 461984
rect 5436 455115 6072 456528
rect 136913 457377 140759 458053
rect 128913 456233 132752 456791
rect 6459 436151 6743 436988
rect 13424 434895 14366 436724
rect 136929 433457 140750 434133
rect 128909 432251 132750 432842
rect 6378 429877 7086 430832
rect 11697 427828 13585 428240
rect 4522 425868 4717 426541
rect 72774 283754 73100 283860
rect 74063 279659 74651 279771
rect 126333 249227 126572 249334
rect 66984 148022 67376 148120
rect 66876 143790 67297 143880
rect 46264 113496 46461 113554
rect 47992 113298 48189 113356
rect 49795 113096 49992 113154
rect 50047 112898 50244 112956
rect 50335 112697 50532 112755
rect 50615 112496 50812 112554
rect 79036 78016 79518 78218
rect 74554 74123 74618 74187
rect 79047 74075 79566 74215
rect 56820 45109 57027 45168
rect 57406 44907 57613 44966
rect 59488 44708 59695 44767
rect 59793 44508 60000 44567
rect 60146 44308 60353 44367
rect 63928 44108 64135 44167
rect 65290 43908 65497 43967
rect 67318 43708 67525 43767
rect 126750 248966 126989 249073
rect 127136 248666 127375 248773
rect 127557 248340 127796 248447
rect 127934 248043 128173 248150
rect 280236 11032 280439 11088
rect 279888 10904 280091 10960
rect 279573 10776 279722 10832
rect 279262 10648 279398 10704
rect 278859 10521 279049 10577
rect 278570 10391 278691 10447
rect 278154 10263 278357 10319
rect 276399 10135 276602 10191
rect 272845 10009 273048 10065
rect 269321 9881 269524 9937
rect 265744 9751 265947 9807
rect 262199 9624 262402 9680
rect 286531 277613 286590 277791
rect 298623 277538 298693 277776
rect 286731 276926 286790 277121
rect 286931 275798 286990 275993
rect 287131 273710 287190 273905
rect 287331 271615 287390 271810
rect 287531 269524 287590 269719
rect 287731 266352 287790 266547
rect 287931 261087 287990 261294
rect 298423 260587 298493 260788
rect 298223 207988 298293 208190
rect 288131 197431 288190 197629
rect 298023 155388 298093 155592
rect 297823 102785 297893 102990
rect 288309 86979 288390 87181
rect 290122 30361 290933 30905
rect 288835 11032 289038 11088
rect 288461 10904 288664 10960
rect 288257 10776 288460 10832
rect 288062 10648 288265 10704
rect 287865 10520 288068 10576
rect 287663 10392 287866 10448
rect 287464 10264 287667 10320
rect 287255 10137 287458 10193
rect 287069 10008 287272 10064
rect 286866 9880 287069 9936
rect 286679 9752 286882 9808
rect 286461 9624 286664 9680
rect 297359 10474 297562 10530
rect 297555 10346 297758 10402
rect 297753 10218 297956 10274
rect 297960 10089 298163 10145
rect 298158 9962 298361 10018
rect 298354 9834 298557 9890
rect 298550 9706 298753 9762
rect 444372 614087 448011 617699
rect 513911 593259 520276 609778
rect 583568 588859 583746 589372
rect 510907 570179 518330 576926
rect 452351 563112 455990 566724
rect 438947 561526 439446 561647
rect 557782 434769 557961 435818
rect 583321 433815 583433 434170
rect 583313 431416 583425 431771
rect 423509 422017 425145 422228
rect 452329 420650 456074 421269
rect 444386 418708 447969 419339
rect 404338 10474 404541 10530
rect 407892 10346 408095 10402
rect 411450 10218 411653 10274
rect 414998 10088 415201 10144
rect 418535 9961 418738 10017
rect 422071 9832 422274 9888
rect 425645 9705 425848 9761
rect 458295 412283 458412 412900
rect 458587 412283 458704 412900
rect 458893 412283 459010 412900
rect 459229 412283 459346 412900
rect 547393 412928 552551 413369
rect 459597 412283 459714 412900
rect 466355 410038 473541 412620
rect 580964 367739 581233 369269
rect 583603 360769 584293 361027
<< metal3 >>
rect 16994 703100 21994 704800
rect 68994 703100 73994 704800
rect 120994 703100 125994 704800
rect 166394 703100 171394 704800
rect 171694 703100 173894 704800
rect 174194 703100 176394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 223394 703100 225594 704800
rect 225894 703100 228094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 325094 703100 327294 704800
rect 327594 703100 329794 704800
rect 330094 703100 335094 704800
rect 414194 703100 419194 704800
rect 466194 703100 471194 704800
rect 18574 687352 19364 703100
rect 71019 691045 71393 703100
rect 71019 690671 117078 691045
rect 18574 686562 105509 687352
rect 800 683312 2500 686042
rect 800 682498 101676 683312
rect 800 681042 2500 682498
rect 800 649314 8531 649442
rect 800 644833 3472 649314
rect 8318 644833 8531 649314
rect 800 644642 8531 644833
rect 800 639260 8531 639442
rect 800 634779 3494 639260
rect 8340 634779 8531 639260
rect 800 634642 8531 634779
rect 800 564868 9296 565042
rect 800 560414 4054 564868
rect 9132 560414 9296 564868
rect 800 560242 9296 560414
rect 800 554880 9296 555042
rect 800 550426 4066 554880
rect 9144 550426 9296 554880
rect 800 550242 9296 550426
rect 800 512330 1280 512442
rect 800 511148 4360 511260
rect 800 509966 1280 510078
rect 800 508784 1280 508896
rect 800 507602 1280 507714
rect 100862 507674 101676 682498
rect 99670 507328 102794 507674
rect 800 506420 1280 506532
rect 99670 504650 100018 507328
rect 102298 504650 102794 507328
rect 99670 504204 102794 504650
rect 28157 492430 38565 492612
rect 28157 486659 28395 492430
rect 38334 486659 38565 492430
rect 28157 486422 38565 486659
rect 18196 479537 18710 479594
rect 18196 478121 18241 479537
rect 18645 478121 18710 479537
rect 18196 478064 18710 478121
rect 4420 475393 12415 475493
rect 4420 470365 6256 475393
rect 12269 470365 12415 475393
rect 4420 470219 12415 470365
rect 18828 475286 24285 475543
rect 18828 470495 19136 475286
rect 24029 470495 24285 475286
rect 18828 470214 24285 470495
rect 15621 469755 15920 469792
rect 838 469256 2512 469278
rect 838 469220 2262 469256
rect 800 469108 2262 469220
rect 838 469013 2262 469108
rect 2247 468578 2262 469013
rect 2494 469013 2512 469256
rect 7459 469236 8334 469270
rect 7459 469100 7494 469236
rect 8300 469220 8334 469236
rect 15621 469220 15660 469755
rect 8300 469108 15660 469220
rect 8300 469100 8334 469108
rect 7459 469073 8334 469100
rect 15621 469083 15660 469108
rect 15889 469083 15920 469755
rect 15621 469053 15920 469083
rect 2494 468578 2511 469013
rect 2247 468557 2511 468578
rect 800 467926 1280 468038
rect 800 466744 1280 466856
rect 800 465562 1280 465674
rect 800 464380 1280 464492
rect 800 463198 1280 463310
rect 7466 461984 8347 462028
rect 7466 461352 7523 461984
rect 8290 461352 8347 461984
rect 7466 461302 8347 461352
rect 5343 456528 6129 456631
rect 5343 455115 5436 456528
rect 6072 455115 6129 456528
rect 5343 455031 6129 455115
rect 43252 452040 45058 452203
rect 43252 443121 43381 452040
rect 44947 443121 45058 452040
rect 104719 448630 105509 686562
rect 103912 448182 106444 448630
rect 103912 446394 104310 448182
rect 106146 446394 106444 448182
rect 103912 446048 106444 446394
rect 6447 436988 6755 437005
rect 6447 436151 6459 436988
rect 6743 436590 6755 436988
rect 13382 436724 14416 436761
rect 6743 436151 12660 436590
rect 6447 436150 12660 436151
rect 6447 436136 6755 436150
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 12220 430688 12660 436150
rect 13382 434895 13424 436724
rect 14366 436708 14416 436724
rect 43252 436708 45058 443121
rect 14366 434902 45058 436708
rect 14366 434895 14416 434902
rect 13382 434848 14416 434895
rect 74070 430688 74510 430689
rect 12220 430248 74510 430688
rect 6302 429814 7162 429877
rect 11637 428240 13660 428297
rect 11637 427828 11697 428240
rect 13585 427828 13660 428240
rect 11637 427782 13660 427828
rect 4484 426541 4759 426575
rect 4484 426125 4522 426541
rect 1061 425998 4522 426125
rect 800 425886 4522 425998
rect 1061 425868 4522 425886
rect 4717 425998 4759 426541
rect 4717 425886 4760 425998
rect 4717 425868 4759 425886
rect 1061 425840 4759 425868
rect 4484 425830 4759 425840
rect 800 424704 1280 424816
rect 800 423522 1280 423634
rect 800 422340 1280 422452
rect 800 421158 1280 421270
rect 800 419976 1280 420088
rect 74070 384820 74510 430248
rect 73769 384777 74673 384820
rect 73769 384033 73831 384777
rect 74622 384033 74673 384777
rect 73769 383978 74673 384033
rect 800 382664 2454 382776
rect 800 381482 1280 381594
rect 800 380300 1280 380412
rect 800 379118 1280 379230
rect 800 377936 1280 378048
rect 800 376754 1280 376866
rect 2342 359856 2454 382664
rect 2342 359756 7556 359856
rect 7456 358678 7556 359756
rect 116704 347944 117078 690671
rect 115878 347766 118262 347944
rect 115878 345626 116072 347766
rect 118072 345626 118262 347766
rect 115878 345460 118262 345626
rect 800 339442 2542 339554
rect 800 338260 1280 338372
rect 800 337078 1280 337190
rect 2341 336449 2542 339442
rect 800 335896 1280 336008
rect 800 334714 1280 334826
rect 800 333532 1280 333644
rect 2342 317188 2542 336449
rect 15656 318928 16056 318962
rect 15656 318190 15702 318928
rect 16022 318190 16056 318928
rect 15656 318140 16056 318190
rect 24316 317188 24516 317838
rect 2342 316988 24516 317188
rect 25156 316348 25356 317838
rect 2342 316148 25356 316348
rect 2342 296332 2578 316148
rect 800 296220 2578 296332
rect 800 295038 1280 295150
rect 800 293856 1280 293968
rect 800 292674 1280 292786
rect 800 291492 1280 291604
rect 800 290310 1280 290422
rect 122792 287156 123728 703100
rect 168369 697685 168783 703100
rect 146740 697271 168783 697685
rect 128832 479922 132832 648476
rect 128832 479271 128886 479922
rect 132750 479271 132832 479922
rect 128832 456791 132832 479271
rect 128832 456233 128913 456791
rect 132752 456233 132832 456791
rect 128832 432842 132832 456233
rect 128832 432251 128909 432842
rect 132750 432251 132832 432842
rect 128832 292274 132832 432251
rect 128832 291646 128946 292274
rect 132748 291646 132832 292274
rect 121856 286830 124852 287156
rect 121856 284192 122182 286830
rect 124562 284192 124852 286830
rect 90434 283976 90842 284006
rect 90434 283872 90462 283976
rect 72760 283860 90462 283872
rect 72760 283754 72774 283860
rect 73100 283754 90462 283860
rect 72760 283742 90462 283754
rect 90434 283662 90462 283742
rect 90814 283662 90842 283976
rect 121856 283880 124852 284192
rect 90434 283634 90842 283662
rect 87789 279902 88281 279936
rect 87789 279785 87851 279902
rect 74040 279771 87851 279785
rect 74040 279659 74063 279771
rect 74651 279659 87851 279771
rect 74040 279641 87851 279659
rect 87789 279549 87851 279641
rect 88235 279549 88281 279902
rect 87789 279501 88281 279549
rect 800 253198 1280 253310
rect 800 252016 1280 252128
rect 800 250834 1280 250946
rect 800 249652 1280 249764
rect 800 248470 1280 248582
rect 52599 248136 52663 251489
rect 55478 248429 55538 251479
rect 55817 248754 55877 251479
rect 56213 249038 56273 251487
rect 60752 249300 60812 251497
rect 126317 249334 126591 249346
rect 126317 249300 126333 249334
rect 60752 249240 126333 249300
rect 126317 249227 126333 249240
rect 126572 249300 126591 249334
rect 126572 249240 128206 249300
rect 126572 249227 126591 249240
rect 126317 249215 126591 249227
rect 126734 249073 127008 249083
rect 126734 249038 126750 249073
rect 56213 248978 126750 249038
rect 126734 248966 126750 248978
rect 126989 249038 127008 249073
rect 126989 248978 128212 249038
rect 126989 248966 127008 248978
rect 126734 248952 127008 248966
rect 127121 248773 127395 248782
rect 127121 248754 127136 248773
rect 55817 248694 127136 248754
rect 127121 248666 127136 248694
rect 127375 248754 127395 248773
rect 127375 248694 128202 248754
rect 127375 248666 127395 248694
rect 127121 248651 127395 248666
rect 127538 248447 127812 248460
rect 127538 248429 127557 248447
rect 55478 248369 127557 248429
rect 127538 248340 127557 248369
rect 127796 248429 127812 248447
rect 127796 248369 128223 248429
rect 127796 248340 127812 248369
rect 127538 248329 127812 248340
rect 127915 248150 128189 248162
rect 127915 248136 127934 248150
rect 52599 248072 127934 248136
rect 127915 248043 127934 248072
rect 128173 248136 128189 248150
rect 128173 248072 128277 248136
rect 128173 248043 128189 248072
rect 127915 248031 128189 248043
rect 800 247288 1280 247400
rect 800 220396 9632 220488
rect 800 215890 4310 220396
rect 9440 215890 9632 220396
rect 800 215688 9632 215890
rect 800 210358 9632 210488
rect 800 205852 4284 210358
rect 9414 205852 9632 210358
rect 800 205688 9632 205852
rect 800 178310 9505 178488
rect 800 173829 3756 178310
rect 8602 173829 9505 178310
rect 800 173688 9505 173829
rect 128832 173511 132832 291646
rect 128832 168834 129023 173511
rect 132621 168834 132832 173511
rect 800 168320 9505 168488
rect 800 163839 3676 168320
rect 8522 163839 9505 168320
rect 800 163688 9505 163839
rect 128832 158446 132832 168834
rect 128832 157840 128914 158446
rect 132770 157840 132832 158446
rect 66970 148120 91441 148132
rect 66970 148022 66984 148120
rect 67376 148022 91441 148120
rect 66970 148010 91441 148022
rect 66865 143880 89792 143889
rect 66865 143790 66876 143880
rect 67297 143790 89792 143880
rect 66865 143780 89792 143790
rect 89683 135800 89792 143780
rect 91319 136400 91441 148010
rect 91130 136386 91694 136400
rect 91130 136206 91146 136386
rect 91678 136206 91694 136386
rect 91130 136192 91694 136206
rect 89683 135780 90361 135800
rect 89683 135626 89701 135780
rect 90336 135626 90361 135780
rect 89683 135606 90361 135626
rect 800 125576 1280 125688
rect 800 124394 1280 124506
rect 800 123212 1280 123324
rect 800 122030 1280 122142
rect 800 120848 1280 120960
rect 800 119666 1280 119778
rect 46323 113564 46387 114487
rect 46257 113554 46470 113564
rect 46257 113496 46264 113554
rect 46461 113496 46470 113554
rect 46257 113489 46470 113496
rect 46323 112434 46387 113489
rect 48059 113364 48123 114487
rect 47985 113356 48198 113364
rect 47985 113298 47992 113356
rect 48189 113298 48198 113356
rect 47985 113289 48198 113298
rect 48059 112434 48123 113289
rect 49863 113164 49923 114487
rect 49788 113154 50001 113164
rect 49788 113096 49795 113154
rect 49992 113096 50001 113154
rect 49788 113089 50001 113096
rect 49863 112434 49923 113089
rect 50111 112964 50171 114487
rect 50040 112956 50253 112964
rect 50040 112898 50047 112956
rect 50244 112898 50253 112956
rect 50040 112889 50253 112898
rect 50111 112434 50171 112889
rect 50395 112764 50455 114487
rect 50326 112755 50539 112764
rect 50326 112697 50335 112755
rect 50532 112697 50539 112755
rect 50326 112689 50539 112697
rect 50395 112434 50455 112689
rect 50677 112564 50737 114487
rect 50608 112554 50821 112564
rect 50608 112496 50615 112554
rect 50812 112496 50821 112554
rect 50608 112489 50821 112496
rect 50677 112434 50737 112489
rect 128832 89424 132832 157840
rect 128832 88794 128928 89424
rect 132734 88794 132832 89424
rect 800 82354 1280 82466
rect 800 81172 1280 81284
rect 800 79990 1280 80102
rect 800 78808 1280 78920
rect 101366 78250 102292 78278
rect 101366 78232 101410 78250
rect 79021 78218 101410 78232
rect 79021 78016 79036 78218
rect 79518 78016 101410 78218
rect 79021 77998 101410 78016
rect 102260 77998 102292 78250
rect 101366 77966 102292 77998
rect 800 77626 1280 77738
rect 800 76444 1280 76556
rect 101158 74261 102354 74287
rect 101158 74230 101199 74261
rect 79030 74215 101199 74230
rect 74549 74187 74623 74192
rect 74549 74123 74554 74187
rect 74618 74123 74623 74187
rect 74549 74118 74623 74123
rect 79030 74075 79047 74215
rect 79566 74075 101199 74215
rect 79030 74060 101199 74075
rect 101158 74009 101199 74060
rect 102314 74009 102354 74261
rect 101158 73980 102354 74009
rect 56877 45175 56937 45901
rect 56808 45168 57039 45175
rect 56808 45109 56820 45168
rect 57027 45109 57039 45168
rect 56808 45099 57039 45109
rect 56877 43671 56937 45099
rect 57470 44975 57534 45905
rect 57397 44966 57628 44975
rect 57397 44907 57406 44966
rect 57613 44907 57628 44966
rect 57397 44899 57628 44907
rect 57470 43671 57534 44899
rect 59553 44775 59613 45901
rect 59479 44767 59710 44775
rect 59479 44708 59488 44767
rect 59695 44708 59710 44767
rect 59479 44699 59710 44708
rect 59553 43671 59613 44699
rect 59861 44575 59921 45901
rect 59782 44567 60013 44575
rect 59782 44508 59793 44567
rect 60000 44508 60013 44567
rect 59782 44499 60013 44508
rect 59861 43671 59921 44499
rect 60211 44375 60271 45901
rect 60135 44367 60366 44375
rect 60135 44308 60146 44367
rect 60353 44308 60366 44367
rect 60135 44299 60366 44308
rect 60211 43671 60271 44299
rect 63998 44175 64058 45910
rect 63917 44167 64148 44175
rect 63917 44108 63928 44167
rect 64135 44108 64148 44167
rect 63917 44099 64148 44108
rect 63998 43671 64058 44099
rect 65358 43975 65418 45905
rect 65278 43967 65509 43975
rect 65278 43908 65290 43967
rect 65497 43908 65509 43967
rect 65278 43899 65509 43908
rect 65358 43671 65418 43899
rect 67398 43775 67458 45910
rect 67309 43767 67540 43775
rect 67309 43708 67318 43767
rect 67525 43708 67540 43767
rect 67309 43699 67540 43708
rect 67398 43671 67458 43699
rect 800 39132 1280 39244
rect 800 37950 1280 38062
rect 800 36768 1280 36880
rect 800 35586 1280 35698
rect 800 34404 1280 34516
rect 128832 34412 132832 88794
rect 136832 644370 140832 645156
rect 136832 639691 136986 644370
rect 140674 639691 140832 644370
rect 136832 481050 140832 639691
rect 136832 480414 136929 481050
rect 140755 480414 140832 481050
rect 136832 458053 140832 480414
rect 136832 457377 136913 458053
rect 140759 457377 140832 458053
rect 136832 434133 140832 457377
rect 136832 433457 136929 434133
rect 140750 433457 140832 434133
rect 136832 362468 140832 433457
rect 144184 384758 145072 384830
rect 144184 384062 144272 384758
rect 144986 384062 145072 384758
rect 144184 383978 145072 384062
rect 136832 361328 136912 362468
rect 140668 361328 140832 362468
rect 136832 293342 140832 361328
rect 136832 292670 136932 293342
rect 140722 292670 140832 293342
rect 136832 159486 140832 292670
rect 136832 158856 136892 159486
rect 140768 158856 140832 159486
rect 136832 90914 140832 158856
rect 144530 136532 144770 383978
rect 146740 146616 147154 697271
rect 220111 693525 220373 703100
rect 160762 693263 220373 693525
rect 160762 277622 161024 693263
rect 331404 680832 331796 703100
rect 415856 686754 416308 703100
rect 467586 686834 468038 703100
rect 511394 698944 516194 704800
rect 511394 693868 511510 698944
rect 516020 693868 516194 698944
rect 511394 693672 516194 693868
rect 521394 698932 526194 704800
rect 567394 703100 572394 704800
rect 521394 693856 521554 698932
rect 526064 693856 526194 698932
rect 521394 693672 526194 693856
rect 415856 686302 427878 686754
rect 331404 680440 424246 680832
rect 423854 607278 424246 680440
rect 422464 606998 426030 607278
rect 422464 604042 422844 606998
rect 425668 604042 426030 606998
rect 422464 603712 426030 604042
rect 427426 510778 427878 686302
rect 430574 686382 468038 686834
rect 426196 510246 429274 510778
rect 426196 507904 426646 510246
rect 428700 507904 429274 510246
rect 426196 507534 429274 507904
rect 284377 478603 284838 478643
rect 284377 477428 284414 478603
rect 284791 477428 284838 478603
rect 284377 477375 284838 477428
rect 164263 299683 283901 300041
rect 160382 277552 161464 277622
rect 160382 276640 160462 277552
rect 161378 276640 161464 277552
rect 160382 276556 161464 276640
rect 145758 146268 148578 146616
rect 145758 143960 146008 146268
rect 148318 143960 148578 146268
rect 145758 143656 148578 143960
rect 144404 136496 144880 136532
rect 144404 136126 144448 136496
rect 144834 136126 144880 136496
rect 144404 136082 144880 136126
rect 136832 90230 136908 90914
rect 140768 90230 140832 90914
rect 136832 34412 140832 90230
rect 144530 78356 144770 136082
rect 144422 78320 144962 78356
rect 144422 77902 144460 78320
rect 144926 77902 144962 78320
rect 144422 77864 144962 77902
rect 144530 77764 144770 77864
rect 160762 66334 161024 276556
rect 164263 274755 164621 299683
rect 165827 297965 283131 298323
rect 164005 274649 164921 274755
rect 164005 273911 164094 274649
rect 164818 273911 164921 274649
rect 164005 273843 164921 273911
rect 165827 136504 166185 297965
rect 165827 135595 165864 136504
rect 166158 135595 166185 136504
rect 165827 135564 166185 135595
rect 166913 296299 282375 296657
rect 166913 74863 167271 296299
rect 280933 295162 281399 295188
rect 280933 293605 280972 295162
rect 281364 293605 281399 295162
rect 280933 293564 281399 293605
rect 280979 267593 281337 293564
rect 282017 270763 282375 296299
rect 282773 272855 283131 297965
rect 283543 274947 283901 299683
rect 284417 276499 284775 477375
rect 430574 430644 431026 686382
rect 467586 686276 468038 686382
rect 568648 683460 569100 703100
rect 433826 683008 569100 683460
rect 429488 430286 432010 430644
rect 429488 428204 429740 430286
rect 431646 428204 432010 430286
rect 429488 427878 432010 428204
rect 423480 422228 425176 422253
rect 423480 422017 423509 422228
rect 425145 422017 425176 422228
rect 423480 421993 425176 422017
rect 423623 387551 423844 421993
rect 285445 387330 423844 387551
rect 285445 276809 285684 387330
rect 433826 376772 434278 683008
rect 583100 680372 584800 683784
rect 436838 679920 584800 680372
rect 432290 376556 435784 376772
rect 432290 373806 432656 376556
rect 435446 373806 435784 376556
rect 432290 373562 435784 373806
rect 436838 287992 437290 679920
rect 583100 678784 584800 679920
rect 573658 645170 584800 645384
rect 444177 640383 448177 641064
rect 573658 640732 573828 645170
rect 578952 640732 584800 645170
rect 573658 640584 584800 640732
rect 444177 635697 444374 640383
rect 448011 635697 448177 640383
rect 444177 617699 448177 635697
rect 444177 614087 444372 617699
rect 448011 614087 448177 617699
rect 438929 561647 439466 561660
rect 438929 561526 438947 561647
rect 439446 561526 439466 561647
rect 438929 561509 439466 561526
rect 438977 384585 439077 561509
rect 444177 419339 448177 614087
rect 444177 418708 444386 419339
rect 447969 418708 448177 419339
rect 438962 384568 439091 384585
rect 438962 384266 438977 384568
rect 439074 384266 439091 384568
rect 438962 384247 439091 384266
rect 435826 287604 440158 287992
rect 435826 284006 436136 287604
rect 439734 284006 440158 287604
rect 435826 283660 440158 284006
rect 285957 277497 286200 279881
rect 286495 277791 288828 277800
rect 286495 277613 286531 277791
rect 286590 277613 288828 277791
rect 297766 277776 298736 277784
rect 297766 277650 298623 277776
rect 286495 277601 288828 277613
rect 298586 277538 298623 277650
rect 298693 277538 298736 277776
rect 298586 277530 298736 277538
rect 285957 277254 288872 277497
rect 297697 277260 298234 277465
rect 298029 277213 298234 277260
rect 286670 277121 288877 277133
rect 286670 276926 286731 277121
rect 286790 276926 288877 277121
rect 298029 277008 299932 277213
rect 286670 276912 288877 276926
rect 285445 276570 288869 276809
rect 284417 276141 288988 276499
rect 286876 275993 288851 276007
rect 286876 275798 286931 275993
rect 286990 275798 288851 275993
rect 286876 275786 288851 275798
rect 283543 274589 288988 274947
rect 287075 273905 288857 273915
rect 287075 273710 287131 273905
rect 287190 273710 288857 273905
rect 287075 273694 288857 273710
rect 282773 272497 288988 272855
rect 287288 271810 288937 271823
rect 287288 271615 287331 271810
rect 287390 271615 288937 271810
rect 287288 271602 288937 271615
rect 282017 270405 288988 270763
rect 287474 269719 288851 269731
rect 287474 269524 287531 269719
rect 287590 269524 288851 269719
rect 287474 269510 288851 269524
rect 280979 267235 288988 267593
rect 287713 266547 288851 266561
rect 287713 266352 287731 266547
rect 287790 266352 288851 266547
rect 287713 266340 288851 266352
rect 284372 261975 288992 262337
rect 297732 261472 299849 261834
rect 287918 261294 288850 261301
rect 287918 261087 287931 261294
rect 287990 261087 288850 261294
rect 287918 261080 288850 261087
rect 297873 260788 298534 260798
rect 297873 260587 298423 260788
rect 298493 260587 298534 260788
rect 297873 260577 298534 260587
rect 297732 208872 299585 209234
rect 297873 208190 298325 208198
rect 297873 207988 298223 208190
rect 298293 207988 298325 208190
rect 297873 207977 298325 207988
rect 284999 198315 288992 198677
rect 288080 197629 288851 197641
rect 288080 197431 288131 197629
rect 288190 197431 288851 197629
rect 288080 197420 288851 197431
rect 297732 156272 299592 156634
rect 297691 155592 298110 155598
rect 297691 155388 298023 155592
rect 298093 155388 298110 155592
rect 297691 155377 298110 155388
rect 297733 103672 299641 104034
rect 285045 87865 288992 88227
rect 288275 87181 288851 87191
rect 288275 86979 288309 87181
rect 288390 86979 288851 87181
rect 288275 86970 288851 86979
rect 166913 73826 166953 74863
rect 167227 73826 167271 74863
rect 166913 73781 167271 73826
rect 159752 66158 162288 66334
rect 159752 63802 159964 66158
rect 162104 63802 162288 66158
rect 159752 63598 162288 63802
rect 285697 46840 289043 47069
rect 297617 46907 301603 47122
rect 444177 34284 448177 418708
rect 452177 566724 456177 637871
rect 573658 635200 584800 635384
rect 573658 630762 573842 635200
rect 578966 630762 584800 635200
rect 573658 630584 584800 630762
rect 513415 609778 520733 610315
rect 513415 593259 513911 609778
rect 520276 593259 520733 609778
rect 513415 592789 520733 593259
rect 584320 590272 584800 590384
rect 583556 589372 583758 589415
rect 583556 588859 583568 589372
rect 583746 589202 583758 589372
rect 583746 589090 584800 589202
rect 583746 588859 583758 589090
rect 583556 588790 583758 588859
rect 584320 587908 584800 588020
rect 584320 586726 584800 586838
rect 584320 585544 584800 585656
rect 584320 584362 584800 584474
rect 510422 576926 518844 577547
rect 510422 570179 510907 576926
rect 518330 570179 518844 576926
rect 510422 569612 518844 570179
rect 452177 563112 452351 566724
rect 455990 563112 456177 566724
rect 452177 421269 456177 563112
rect 549766 558443 549932 573064
rect 452177 420650 452329 421269
rect 456074 420650 456177 421269
rect 452177 191899 456177 420650
rect 458275 558277 549932 558443
rect 458275 412900 458441 558277
rect 550058 558151 550224 573064
rect 458275 412283 458295 412900
rect 458412 412283 458441 412900
rect 458275 412236 458441 412283
rect 458567 557985 550224 558151
rect 458567 412900 458733 557985
rect 550363 557846 550529 573064
rect 458567 412283 458587 412900
rect 458704 412283 458733 412900
rect 458567 412236 458733 412283
rect 458872 557680 550529 557846
rect 458872 412900 459038 557680
rect 550698 557511 550864 573064
rect 458872 412283 458893 412900
rect 459010 412283 459038 412900
rect 458872 412236 459038 412283
rect 459207 557345 550864 557511
rect 459207 412900 459373 557345
rect 552764 557145 552972 573064
rect 459207 412283 459229 412900
rect 459346 412283 459373 412900
rect 459207 412236 459373 412283
rect 459573 556937 552972 557145
rect 459573 412900 459781 556937
rect 575498 556038 584800 556162
rect 575498 551600 575644 556038
rect 580768 551600 584800 556038
rect 575498 551362 584800 551600
rect 575498 546004 584800 546162
rect 575498 541566 575630 546004
rect 580754 541566 584800 546004
rect 575498 541362 584800 541566
rect 584320 500850 584800 500962
rect 557755 499780 584508 499829
rect 557755 499668 584800 499780
rect 557755 499598 584508 499668
rect 557755 435818 557986 499598
rect 584320 498486 584800 498598
rect 584320 497304 584800 497416
rect 584320 496122 584800 496234
rect 584320 494940 584800 495052
rect 584320 456428 584800 456540
rect 584320 455246 584800 455358
rect 584320 454064 584800 454176
rect 584320 452882 584800 452994
rect 557755 434769 557782 435818
rect 557961 434769 557986 435818
rect 557755 434744 557986 434769
rect 583321 451700 584800 451812
rect 475894 434151 479604 434328
rect 583321 434178 583433 451700
rect 584320 450518 584800 450630
rect 475894 425383 476138 434151
rect 479384 425383 479604 434151
rect 583313 434170 583443 434178
rect 583313 433815 583321 434170
rect 583433 433815 583443 434170
rect 583313 433801 583443 433815
rect 583321 433794 583433 433801
rect 583313 431779 583425 431796
rect 583305 431771 583434 431779
rect 583305 431416 583313 431771
rect 583425 431416 583434 431771
rect 583305 431407 583434 431416
rect 475894 425155 479604 425383
rect 475901 413650 478420 425155
rect 475901 413369 552664 413650
rect 475901 412928 547393 413369
rect 552551 412928 552664 413369
rect 475901 412913 552664 412928
rect 459573 412283 459597 412900
rect 459714 412283 459781 412900
rect 459573 412236 459781 412283
rect 466206 412620 473703 412769
rect 466206 410038 466355 412620
rect 473541 410038 473703 412620
rect 466206 409865 473703 410038
rect 583313 407390 583425 431407
rect 584320 412006 584800 412118
rect 584320 410824 584800 410936
rect 584320 409642 584800 409754
rect 584320 408460 584800 408572
rect 583313 407278 584800 407390
rect 584320 406096 584800 406208
rect 580563 384575 581315 384602
rect 580563 384268 580603 384575
rect 581287 384268 581315 384575
rect 580563 384240 581315 384268
rect 580951 369297 581251 384240
rect 580930 369269 581274 369297
rect 580930 367739 580964 369269
rect 581233 367739 581274 369269
rect 580930 367703 581274 367739
rect 584320 365584 584800 365696
rect 584320 364402 584800 364514
rect 584320 363220 584800 363332
rect 584320 362038 584800 362150
rect 583575 361027 584320 361051
rect 583575 360769 583603 361027
rect 584293 360968 584320 361027
rect 584293 360856 584800 360968
rect 584293 360769 584320 360856
rect 583575 360746 584320 360769
rect 584320 359674 584800 359786
rect 573750 326498 582242 326852
rect 581888 315867 582242 326498
rect 584320 320362 584800 320474
rect 584320 319180 584800 319292
rect 584320 317998 584800 318110
rect 584320 316816 584800 316928
rect 581888 315746 584383 315867
rect 581888 315634 584800 315746
rect 581888 315513 584383 315634
rect 584320 314452 584800 314564
rect 584320 275940 584800 276052
rect 584320 274758 584800 274870
rect 584320 273576 584800 273688
rect 584320 272394 584800 272506
rect 584320 271212 584800 271324
rect 584320 270030 584800 270142
rect 574794 240690 584800 240830
rect 574794 236252 574934 240690
rect 580058 236252 584800 240690
rect 574794 236030 584800 236252
rect 574794 230660 584800 230830
rect 574794 226222 574962 230660
rect 580086 226222 584800 230660
rect 574794 226030 584800 226222
rect 574794 196850 584800 197030
rect 574794 192412 574896 196850
rect 580020 192412 584800 196850
rect 574794 192230 584800 192412
rect 452177 187251 452333 191899
rect 455990 187251 456177 191899
rect 452177 34284 456177 187251
rect 574794 186806 584800 187030
rect 574794 182368 574908 186806
rect 580032 182368 584800 186806
rect 574794 182230 584800 182368
rect 574794 152256 584800 152430
rect 574794 147818 575156 152256
rect 580280 147818 584800 152256
rect 574794 147630 584800 147818
rect 574794 142194 584800 142430
rect 574794 137756 575102 142194
rect 580226 137756 584800 142194
rect 574794 137630 584800 137756
rect 584320 95918 584800 96030
rect 584320 94736 584800 94848
rect 584320 93554 584800 93666
rect 584320 92372 584800 92484
rect 584320 51260 584800 51372
rect 584320 50078 584800 50190
rect 584320 48896 584800 49008
rect 584320 47714 584800 47826
rect 800 33222 1280 33334
rect 290073 30905 290992 30949
rect 290073 30361 290122 30905
rect 290933 30682 290992 30905
rect 290933 30361 290994 30682
rect 290073 30317 290994 30361
rect 2528 18157 3384 18189
rect 2528 17976 2562 18157
rect 1114 17822 2562 17976
rect 800 17710 2562 17822
rect 1114 17563 2562 17710
rect 2528 17264 2562 17563
rect 3344 17264 3384 18157
rect 2528 17233 3384 17264
rect 290074 18165 290994 30317
rect 584320 24802 584800 24914
rect 584320 23620 584800 23732
rect 584320 22438 584800 22550
rect 584320 21256 584800 21368
rect 584320 20074 584800 20186
rect 584320 18892 584800 19004
rect 290074 17259 290103 18165
rect 290967 17259 290994 18165
rect 584320 17710 584800 17822
rect 290074 17234 290994 17259
rect 800 16528 1280 16640
rect 584320 16528 584800 16640
rect 800 15346 1280 15458
rect 584320 15346 584800 15458
rect 800 14164 1280 14276
rect 584320 14164 584800 14276
rect 800 12982 1280 13094
rect 584320 12982 584800 13094
rect 800 11800 1280 11912
rect 584320 11800 584800 11912
rect 280227 11091 280448 11093
rect 288826 11091 289047 11093
rect 262134 11088 289047 11091
rect 262134 11032 280236 11088
rect 280439 11032 288835 11088
rect 289038 11032 289047 11088
rect 262134 11027 289047 11032
rect 279879 10963 280100 10965
rect 288452 10963 288673 10965
rect 262134 10960 288997 10963
rect 262134 10904 279888 10960
rect 280091 10904 288461 10960
rect 288664 10904 288997 10960
rect 262134 10899 288997 10904
rect 279510 10835 279731 10837
rect 288248 10835 288469 10837
rect 262134 10832 288997 10835
rect 262134 10776 279573 10832
rect 279722 10776 288257 10832
rect 288460 10776 288997 10832
rect 262134 10771 288997 10776
rect 800 10618 1280 10730
rect 279186 10707 279407 10709
rect 288053 10707 288274 10709
rect 262134 10704 288997 10707
rect 262134 10648 279262 10704
rect 279398 10648 288062 10704
rect 288265 10648 288997 10704
rect 262134 10643 288997 10648
rect 584320 10618 584800 10730
rect 278837 10579 279058 10582
rect 287856 10579 288077 10581
rect 262134 10577 288997 10579
rect 262134 10521 278859 10577
rect 279049 10576 288997 10577
rect 279049 10521 287865 10576
rect 262134 10520 287865 10521
rect 288068 10520 288997 10576
rect 297350 10532 297571 10535
rect 404329 10532 404550 10535
rect 262134 10515 288997 10520
rect 297282 10530 425861 10532
rect 297282 10474 297359 10530
rect 297562 10474 404338 10530
rect 404541 10474 425861 10530
rect 297282 10468 425861 10474
rect 278479 10451 278700 10452
rect 287654 10451 287875 10453
rect 262134 10448 288997 10451
rect 262134 10447 287663 10448
rect 262134 10391 278570 10447
rect 278691 10392 287663 10447
rect 287866 10392 288997 10448
rect 297546 10404 297767 10407
rect 407883 10404 408104 10407
rect 278691 10391 288997 10392
rect 262134 10387 288997 10391
rect 297282 10402 425861 10404
rect 278479 10386 278700 10387
rect 297282 10346 297555 10402
rect 297758 10346 407892 10402
rect 408095 10346 425861 10402
rect 297282 10340 425861 10346
rect 278145 10323 278366 10324
rect 287455 10323 287676 10325
rect 262134 10320 288997 10323
rect 262134 10319 287464 10320
rect 262134 10263 278154 10319
rect 278357 10264 287464 10319
rect 287667 10264 288997 10320
rect 297744 10276 297965 10279
rect 411441 10276 411662 10279
rect 278357 10263 288997 10264
rect 262134 10259 288997 10263
rect 297282 10274 425861 10276
rect 278145 10258 278366 10259
rect 297282 10218 297753 10274
rect 297956 10218 411450 10274
rect 411653 10218 425861 10274
rect 297282 10212 425861 10218
rect 276390 10195 276611 10196
rect 287246 10195 287467 10198
rect 262134 10193 288997 10195
rect 262134 10191 287255 10193
rect 262134 10135 276399 10191
rect 276602 10137 287255 10191
rect 287458 10137 288997 10193
rect 297951 10148 298172 10150
rect 414989 10148 415210 10149
rect 276602 10135 288997 10137
rect 262134 10131 288997 10135
rect 297282 10145 425861 10148
rect 276390 10130 276611 10131
rect 297282 10089 297960 10145
rect 298163 10144 425861 10145
rect 298163 10089 414998 10144
rect 297282 10088 414998 10089
rect 415201 10088 425861 10144
rect 297282 10084 425861 10088
rect 414989 10083 415210 10084
rect 272836 10067 273050 10070
rect 287060 10067 287281 10069
rect 262134 10065 288997 10067
rect 262134 10009 272845 10065
rect 273048 10064 288997 10065
rect 273048 10009 287069 10064
rect 262134 10008 287069 10009
rect 287272 10008 288997 10064
rect 298149 10020 298370 10023
rect 418526 10020 418747 10022
rect 262134 10003 288997 10008
rect 297282 10018 425861 10020
rect 297282 9962 298158 10018
rect 298361 10017 425861 10018
rect 298361 9962 418535 10017
rect 297282 9961 418535 9962
rect 418738 9961 425861 10017
rect 297282 9956 425861 9961
rect 269312 9939 269533 9942
rect 286857 9939 287078 9941
rect 262134 9937 288997 9939
rect 262134 9881 269321 9937
rect 269524 9936 288997 9937
rect 269524 9881 286866 9936
rect 262134 9880 286866 9881
rect 287069 9880 288997 9936
rect 298345 9892 298566 9895
rect 422062 9892 422283 9893
rect 262134 9875 288997 9880
rect 297282 9890 425861 9892
rect 297282 9834 298354 9890
rect 298557 9888 425861 9890
rect 298557 9834 422071 9888
rect 297282 9832 422071 9834
rect 422274 9832 425861 9888
rect 297282 9828 425861 9832
rect 422062 9827 422283 9828
rect 265735 9811 265956 9812
rect 286670 9811 286891 9813
rect 262134 9808 288997 9811
rect 262134 9807 286679 9808
rect 262134 9751 265744 9807
rect 265947 9752 286679 9807
rect 286882 9752 288997 9808
rect 298541 9764 298762 9767
rect 425636 9764 425857 9766
rect 265947 9751 288997 9752
rect 262134 9747 288997 9751
rect 297282 9762 425861 9764
rect 265735 9746 265956 9747
rect 297282 9706 298550 9762
rect 298753 9761 425861 9762
rect 298753 9706 425645 9761
rect 297282 9705 425645 9706
rect 425848 9705 425861 9761
rect 297282 9700 425861 9705
rect 262190 9683 262411 9685
rect 286452 9683 286673 9685
rect 262134 9680 288997 9683
rect 262134 9624 262199 9680
rect 262402 9624 286461 9680
rect 286664 9624 288997 9680
rect 262134 9619 288997 9624
rect 800 9436 1280 9548
rect 584320 9436 584800 9548
rect 800 8254 1280 8366
rect 584320 8254 584800 8366
rect 800 7072 1280 7184
rect 584320 7072 584800 7184
rect 800 5890 1280 6002
rect 584320 5890 584800 6002
rect 800 4708 1280 4820
rect 584320 4708 584800 4820
rect 800 3526 1280 3638
rect 584320 3526 584800 3638
rect 800 2344 1280 2456
rect 584320 2344 584800 2456
<< via3 >>
rect 3472 644833 8318 649314
rect 3494 634779 8340 639260
rect 4054 560414 9132 564868
rect 4066 550426 9144 554880
rect 100018 504650 102298 507328
rect 28395 486659 38334 492430
rect 18241 478121 18645 479537
rect 6256 470365 12269 475393
rect 19136 470495 24029 475286
rect 7523 461352 8290 461984
rect 5436 455115 6072 456528
rect 43381 443121 44947 452040
rect 104310 446394 106146 448182
rect 6378 429877 7086 430832
rect 11697 427828 13585 428240
rect 73831 384033 74622 384777
rect 116072 345626 118072 347766
rect 15702 318190 16022 318928
rect 128946 291646 132748 292274
rect 122182 284192 124562 286830
rect 90462 283662 90814 283976
rect 87851 279549 88235 279902
rect 4310 215890 9440 220396
rect 4284 205852 9414 210358
rect 3756 173829 8602 178310
rect 129023 168834 132621 173511
rect 3676 163839 8522 168320
rect 128914 157840 132770 158446
rect 91146 136206 91678 136386
rect 89701 135626 90336 135780
rect 128928 88794 132734 89424
rect 101410 77998 102260 78250
rect 101199 74009 102314 74261
rect 136986 639691 140674 644370
rect 144272 384062 144986 384758
rect 136912 361328 140668 362468
rect 136932 292670 140722 293342
rect 136892 158856 140768 159486
rect 511510 693868 516020 698944
rect 521554 693856 526064 698932
rect 422844 604042 425668 606998
rect 426646 507904 428700 510246
rect 284414 477428 284791 478603
rect 160462 276640 161378 277552
rect 146008 143960 148318 146268
rect 144448 136126 144834 136496
rect 136908 90230 140768 90914
rect 144460 77902 144926 78320
rect 164094 273911 164818 274649
rect 165864 135595 166158 136504
rect 280972 293605 281364 295162
rect 429740 428204 431646 430286
rect 432656 373806 435446 376556
rect 573828 640732 578952 645170
rect 444374 635697 448011 640383
rect 438977 384266 439074 384568
rect 436136 284006 439734 287604
rect 166953 73826 167227 74863
rect 159964 63802 162104 66158
rect 573842 630762 578966 635200
rect 513911 593259 520276 609778
rect 510907 570179 518330 576926
rect 575644 551600 580768 556038
rect 575630 541566 580754 546004
rect 476138 425383 479384 434151
rect 466355 410038 473541 412620
rect 580603 384268 581287 384575
rect 574934 236252 580058 240690
rect 574962 226222 580086 230660
rect 574896 192412 580020 196850
rect 452333 187251 455990 191899
rect 574908 182368 580032 186806
rect 575156 147818 580280 152256
rect 575102 137756 580226 142194
rect 2562 17264 3344 18157
rect 290103 17259 290967 18165
<< metal4 >>
rect 166394 703100 171394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 330094 703100 335094 704800
rect 511354 698944 526180 699076
rect 511354 693868 511510 698944
rect 516020 698932 526180 698944
rect 516020 693868 516456 698932
rect 511354 693856 516456 693868
rect 520966 693856 521554 698932
rect 526064 693856 526180 698932
rect 511354 693672 526180 693856
rect 3308 649314 8544 649486
rect 3308 644833 3472 649314
rect 8318 644833 8544 649314
rect 3308 644534 8544 644833
rect 573700 645170 579138 645386
rect 3308 644370 141468 644534
rect 3308 639691 136986 644370
rect 140674 639691 141468 644370
rect 573700 640732 573828 645170
rect 578952 640732 579138 645170
rect 573700 640538 579138 640732
rect 3308 639534 141468 639691
rect 443754 640383 579138 640538
rect 3308 639260 8544 639534
rect 3308 634779 3494 639260
rect 8340 634779 8544 639260
rect 443754 635697 444374 640383
rect 448011 635697 579138 640383
rect 443754 635538 579138 635697
rect 3308 634618 8544 634779
rect 573700 635200 579138 635538
rect 573700 630762 573842 635200
rect 578966 630762 579138 635200
rect 573700 630566 579138 630762
rect 97611 601186 169654 610368
rect 417050 610315 515494 610324
rect 417050 609778 520733 610315
rect 417050 606998 513911 609778
rect 417050 604042 422844 606998
rect 425668 604042 513911 606998
rect 417050 601142 513911 604042
rect 513415 593259 513911 601142
rect 520276 593259 520733 609778
rect 513415 592789 520733 593259
rect 466103 577278 518844 577547
rect 466103 569837 466468 577278
rect 473449 576926 518844 577278
rect 473449 570179 510907 576926
rect 518330 570179 518844 576926
rect 473449 569837 518844 570179
rect 466103 569612 518844 569837
rect 3906 564868 9344 565044
rect 3906 560414 4054 564868
rect 9132 560414 9344 564868
rect 3906 560048 9344 560414
rect 3906 555362 4066 560048
rect 9170 555362 9344 560048
rect 3906 554880 9344 555362
rect 3906 550426 4066 554880
rect 9144 550426 9344 554880
rect 3906 550224 9344 550426
rect 466125 560021 473749 560331
rect 466125 553646 466599 560021
rect 473439 553646 473749 560021
rect 466125 530621 473749 553646
rect 575502 556038 580940 556170
rect 575502 551600 575644 556038
rect 580768 551600 580940 556038
rect 575502 550970 580940 551600
rect 575502 546532 575622 550970
rect 580746 546532 580940 550970
rect 575502 546004 580940 546532
rect 575502 541566 575630 546004
rect 580754 541566 580940 546004
rect 575502 541350 580940 541566
rect 466125 523885 466547 530621
rect 473413 523885 473749 530621
rect 466125 523522 473749 523885
rect 60811 507328 169654 510368
rect 60811 504650 100018 507328
rect 102298 504650 169654 507328
rect 417050 510246 486115 514324
rect 417050 507904 426646 510246
rect 428700 507904 486115 510246
rect 417050 505142 486115 507904
rect 60811 501186 169654 504650
rect 60811 494403 69993 501186
rect 27578 492430 69993 494403
rect 27578 486659 28395 492430
rect 38334 486659 69993 492430
rect 27578 485221 69993 486659
rect 18196 479537 18710 479594
rect 18196 478121 18241 479537
rect 18645 478497 18710 479537
rect 284377 478603 284838 478643
rect 284377 478497 284414 478603
rect 18645 478121 284414 478497
rect 18196 478067 284414 478121
rect 18196 478064 18710 478067
rect 284377 477428 284414 478067
rect 284791 477428 284838 478603
rect 284377 477375 284838 477428
rect 4420 475393 114425 475493
rect 4420 470365 6256 475393
rect 12269 475380 114425 475393
rect 12269 475286 106611 475380
rect 12269 470495 19136 475286
rect 24029 470495 106611 475286
rect 12269 470365 106611 470495
rect 4420 470309 106611 470365
rect 113894 470309 114425 475380
rect 4420 470219 114425 470309
rect 150797 462824 158032 462940
rect 150797 462028 150899 462824
rect 7466 461984 150899 462028
rect 7466 461352 7523 461984
rect 8290 461395 150899 461984
rect 157916 462028 158032 462824
rect 157916 461395 158180 462028
rect 8290 461352 158180 461395
rect 7466 461302 158180 461352
rect 150797 461301 158032 461302
rect 5343 456528 6129 456631
rect 5343 455115 5436 456528
rect 6072 455757 6129 456528
rect 106510 455757 114021 455761
rect 6072 455661 114021 455757
rect 6072 455115 106619 455661
rect 5343 455031 106619 455115
rect 106510 454319 106619 455031
rect 113903 454319 114021 455661
rect 106510 454196 114021 454319
rect 42751 452040 169654 452168
rect 42751 443121 43381 452040
rect 44947 448182 169654 452040
rect 44947 446394 104310 448182
rect 106146 446394 169654 448182
rect 44947 443121 169654 446394
rect 42751 442986 169654 443121
rect 106528 441575 114020 441685
rect 106528 440841 106630 441575
rect 81054 440408 106630 440841
rect 113902 440841 114020 441575
rect 113902 440408 114120 440841
rect 81054 440326 114120 440408
rect 150780 440395 158029 440524
rect 6302 430832 7162 430887
rect 6302 429877 6378 430832
rect 7086 429877 7162 430832
rect 6302 429814 7162 429877
rect 6469 427411 7004 429814
rect 81054 428297 81569 440326
rect 106528 440321 114020 440326
rect 150780 439439 150941 440395
rect 11637 428240 81569 428297
rect 11637 427828 11697 428240
rect 13585 427828 81569 428240
rect 11637 427782 81569 427828
rect 82329 439040 150941 439439
rect 157881 439040 158029 440395
rect 82329 438906 158029 439040
rect 82329 438904 157979 438906
rect 82329 427411 82864 438904
rect 6469 426876 82864 427411
rect 417050 434151 479733 434324
rect 417050 430286 476138 434151
rect 417050 428204 429740 430286
rect 431646 428204 476138 430286
rect 417050 425383 476138 428204
rect 479384 425383 479733 434151
rect 417050 425142 479733 425383
rect 466206 412620 473703 412769
rect 466206 410038 466355 412620
rect 473541 410038 473703 412620
rect 466206 409865 473703 410038
rect 73769 384777 74673 384820
rect 73769 384033 73831 384777
rect 74622 384569 74673 384777
rect 144184 384758 145072 384830
rect 144184 384569 144272 384758
rect 74622 384262 144272 384569
rect 74622 384033 74673 384262
rect 73769 383978 74673 384033
rect 144184 384062 144272 384262
rect 144986 384569 145072 384758
rect 438962 384569 439091 384585
rect 580563 384575 581315 384602
rect 580563 384569 580603 384575
rect 144986 384568 580603 384569
rect 144986 384266 438977 384568
rect 439074 384268 580603 384568
rect 581287 384268 581315 384575
rect 439074 384266 581315 384268
rect 144986 384262 581315 384266
rect 144986 384062 145072 384262
rect 438962 384247 439091 384262
rect 580563 384240 581315 384262
rect 144184 383978 145072 384062
rect 417050 376556 485757 380324
rect 417050 373806 432656 376556
rect 435446 373806 485757 376556
rect 417050 371142 485757 373806
rect 5812 362468 140772 362536
rect 5812 361328 136912 362468
rect 140668 361328 140772 362468
rect 5812 361280 140772 361328
rect 5816 358120 6116 361280
rect 55959 350620 169654 352368
rect 51456 350180 169654 350620
rect 55959 347766 169654 350180
rect 55959 345626 116072 347766
rect 118072 345626 169654 347766
rect 55959 343186 169654 345626
rect 6486 313656 7274 319328
rect 15657 318928 16052 319021
rect 15657 318190 15702 318928
rect 16022 318190 16052 318928
rect 15657 315893 16052 318190
rect 15657 315498 126297 315893
rect 6486 313538 114161 313656
rect 6486 310456 106704 313538
rect 113848 310456 114161 313538
rect 6486 310314 114161 310456
rect 67876 295916 118290 296316
rect 69687 295456 117584 295856
rect 69687 294996 93810 295396
rect 69687 294536 92294 294936
rect 90434 283976 90842 284006
rect 90434 283662 90462 283976
rect 90814 283662 90842 283976
rect 90434 283634 90842 283662
rect 87789 279902 88281 279936
rect 87789 279549 87851 279902
rect 88235 279549 88281 279902
rect 87789 279501 88281 279549
rect 87936 274383 88155 279501
rect 90582 277122 90718 283634
rect 91894 279548 92294 294536
rect 93410 290368 93810 294996
rect 117184 292132 117584 295456
rect 117890 293226 118290 295916
rect 125902 295188 126297 315498
rect 322545 298063 326987 298248
rect 322545 297074 322730 298063
rect 125902 295162 281399 295188
rect 125902 294793 280972 295162
rect 280933 293605 280972 294793
rect 281364 293605 281399 295162
rect 280933 293564 281399 293605
rect 291775 294833 322730 297074
rect 136836 293342 140832 293416
rect 136836 293226 136932 293342
rect 117890 292826 136932 293226
rect 136836 292670 136932 292826
rect 140722 292670 140832 293342
rect 136836 292568 140832 292670
rect 128830 292274 132834 292366
rect 128830 292132 128946 292274
rect 117184 291732 128946 292132
rect 128830 291646 128946 291732
rect 132748 291646 132834 292274
rect 128830 291560 132834 291646
rect 93325 286830 169654 290368
rect 93325 284192 122182 286830
rect 124562 284192 169654 286830
rect 93325 281186 169654 284192
rect 106532 280018 114000 280088
rect 106532 279548 106628 280018
rect 91894 279148 106628 279548
rect 106532 278712 106628 279148
rect 113928 278712 114000 280018
rect 106532 278628 114000 278712
rect 291775 278473 293460 294833
rect 322545 293627 322730 294833
rect 326798 293627 326987 298063
rect 322545 293467 326987 293627
rect 417050 287604 481818 290324
rect 417050 284006 436136 287604
rect 439734 284006 481818 287604
rect 293611 281232 313097 281381
rect 293611 279800 306274 281232
rect 312971 279800 313097 281232
rect 417050 281142 481818 284006
rect 293611 279696 313097 279800
rect 293611 278473 295296 279696
rect 160382 277552 161464 277622
rect 160382 277122 160462 277552
rect 90582 276986 160462 277122
rect 160382 276640 160462 276986
rect 161378 276640 161464 277552
rect 160382 276556 161464 276640
rect 164005 274649 164921 274755
rect 164005 274383 164094 274649
rect 87936 274164 164094 274383
rect 164005 273911 164094 274164
rect 164818 273911 164921 274649
rect 164005 273843 164921 273911
rect 466249 255107 473735 255449
rect 466249 247031 466498 255107
rect 473424 247031 473735 255107
rect 106501 232157 114025 232502
rect 106501 224846 106878 232157
rect 113676 224846 114025 232157
rect 4152 220396 9590 220510
rect 4152 215890 4310 220396
rect 9440 215890 9590 220396
rect 4152 215436 9590 215890
rect 4152 210800 4232 215436
rect 9414 210800 9590 215436
rect 4152 210358 9590 210800
rect 4152 205852 4284 210358
rect 9414 205852 9590 210358
rect 4152 205690 9590 205852
rect 106501 201306 114025 224846
rect 466249 221314 473735 247031
rect 574774 240690 580212 240866
rect 574774 236252 574934 240690
rect 580058 236252 580212 240690
rect 574774 235522 580212 236252
rect 574774 231084 574962 235522
rect 580086 231084 580212 235522
rect 574774 230660 580212 231084
rect 574774 226222 574962 230660
rect 580086 226222 580212 230660
rect 574774 226046 580212 226222
rect 466249 211313 466529 221314
rect 473424 211313 473735 221314
rect 466249 210816 473735 211313
rect 106501 194909 106922 201306
rect 113632 194909 114025 201306
rect 106501 194569 114025 194909
rect 574748 196850 580186 197028
rect 574748 192412 574896 196850
rect 580020 192412 580186 196850
rect 574748 192076 580186 192412
rect 451946 191899 580186 192076
rect 451946 187251 452333 191899
rect 455990 187251 580186 191899
rect 451946 187076 580186 187251
rect 574748 186806 580186 187076
rect 574748 182368 574908 186806
rect 580032 182368 580186 186806
rect 574748 182208 580186 182368
rect 3532 178310 8768 178430
rect 3532 173829 3756 178310
rect 8602 173829 8768 178310
rect 3532 173694 8768 173829
rect 3532 173511 133180 173694
rect 3532 168834 129023 173511
rect 132621 168834 133180 173511
rect 3532 168694 133180 168834
rect 3532 168320 8768 168694
rect 3532 163839 3676 168320
rect 8522 163839 8768 168320
rect 3532 163716 8768 163839
rect 417050 161142 483967 170324
rect 136834 159486 140834 159536
rect 136834 159359 136892 159486
rect 60888 158959 136892 159359
rect 62646 158499 123632 158899
rect 136834 158856 136892 158959
rect 140768 158856 140834 159486
rect 136834 158788 140834 158856
rect 62656 158039 94968 158439
rect 62656 157579 93408 157979
rect 93008 138968 93408 157579
rect 94568 150368 94968 158039
rect 123232 158340 123632 158499
rect 128830 158446 132832 158498
rect 128830 158340 128914 158446
rect 123232 157940 128914 158340
rect 128830 157840 128914 157940
rect 132770 157840 132832 158446
rect 128830 157786 132832 157840
rect 574794 152256 580634 152400
rect 94396 146268 169654 150368
rect 94396 143960 146008 146268
rect 148318 143960 169654 146268
rect 94396 141186 169654 143960
rect 574794 147818 575156 152256
rect 580280 147818 580634 152256
rect 574794 147254 580634 147818
rect 574794 142816 575132 147254
rect 580256 142816 580634 147254
rect 574794 142194 580634 142816
rect 106506 139242 114044 139300
rect 106506 138968 106578 139242
rect 93008 138568 106578 138968
rect 106506 138416 106578 138568
rect 113928 138416 114044 139242
rect 106506 138340 114044 138416
rect 574794 137756 575102 142194
rect 580226 137756 580634 142194
rect 574794 137630 580634 137756
rect 144404 136496 144880 136532
rect 144404 136400 144448 136496
rect 91130 136386 144448 136400
rect 91130 136206 91146 136386
rect 91678 136206 144448 136386
rect 91130 136192 144448 136206
rect 144404 136126 144448 136192
rect 144834 136126 144880 136496
rect 144404 136082 144880 136126
rect 165828 136504 166185 136533
rect 89683 135791 90361 135800
rect 165828 135791 165864 136504
rect 89683 135780 165864 135791
rect 89683 135626 89701 135780
rect 90336 135637 165864 135780
rect 90336 135626 90361 135637
rect 89683 135606 90361 135626
rect 165828 135595 165864 135637
rect 166158 135595 166185 136504
rect 165828 135565 166185 135595
rect 136824 90914 140862 90990
rect 136824 90738 136908 90914
rect 72886 90338 136908 90738
rect 74623 89878 126258 90278
rect 136824 90230 136908 90338
rect 140768 90738 140862 90914
rect 140768 90338 140868 90738
rect 140768 90230 140862 90338
rect 136824 90146 140862 90230
rect 74623 89418 95760 89818
rect 74623 88958 93058 89358
rect 92658 59020 93058 88958
rect 95360 70368 95760 89418
rect 125858 89290 126258 89878
rect 128830 89424 132828 89500
rect 128830 89290 128928 89424
rect 125858 88890 128928 89290
rect 128830 88794 128928 88890
rect 132734 88794 132828 89424
rect 128830 88718 132828 88794
rect 144422 78320 144962 78356
rect 144422 78280 144460 78320
rect 101366 78250 144460 78280
rect 101366 77998 101410 78250
rect 102260 77998 144460 78250
rect 101366 77966 144460 77998
rect 144422 77902 144460 77966
rect 144926 77902 144962 78320
rect 144422 77864 144962 77902
rect 166912 74863 167279 74900
rect 101158 74261 102354 74287
rect 101158 74009 101199 74261
rect 102314 74236 102354 74261
rect 166912 74236 166953 74863
rect 102314 74036 166953 74236
rect 102314 74009 102354 74036
rect 101158 73980 102354 74009
rect 166912 73826 166953 74036
rect 167227 73826 167279 74863
rect 166912 73780 167279 73826
rect 95111 66158 169654 70368
rect 95111 63802 159964 66158
rect 162104 63802 169654 66158
rect 95111 61186 169654 63802
rect 417050 61142 529090 70324
rect 106524 59276 114056 59366
rect 106524 59020 106648 59276
rect 92658 58620 106648 59020
rect 106524 58454 106648 58620
rect 113876 58454 114056 59276
rect 106524 58360 114056 58454
rect 426799 39173 434047 39338
rect 291775 24480 293460 32589
rect 293611 27790 295296 32589
rect 426799 32240 426979 39173
rect 433851 32240 434047 39173
rect 426799 32090 434047 32240
rect 293611 27651 313157 27790
rect 293611 26209 306753 27651
rect 313014 26209 313157 27651
rect 293611 26105 313157 26209
rect 428910 24480 430595 32090
rect 291775 22795 430595 24480
rect 2527 18165 291000 18190
rect 2527 18157 290103 18165
rect 2527 17264 2562 18157
rect 3344 17264 290103 18157
rect 2527 17259 290103 17264
rect 290967 17259 291000 18165
rect 2527 17232 291000 17259
<< via4 >>
rect 516456 693856 520966 698932
rect 466468 569837 473449 577278
rect 4066 555362 9170 560048
rect 466599 553646 473439 560021
rect 575622 546532 580746 550970
rect 466547 523885 473413 530621
rect 106611 470309 113894 475380
rect 150899 461395 157916 462824
rect 106619 454319 113903 455661
rect 106630 440408 113902 441575
rect 150941 439040 157881 440395
rect 466355 410038 473541 412620
rect 106704 310456 113848 313538
rect 106628 278712 113928 280018
rect 322730 293627 326798 298063
rect 306274 279800 312971 281232
rect 466498 247031 473424 255107
rect 106878 224846 113676 232157
rect 4232 210800 9414 215436
rect 574962 231084 580086 235522
rect 466529 211313 473424 221314
rect 106922 194909 113632 201306
rect 575132 142816 580256 147254
rect 106578 138416 113928 139242
rect 106648 58454 113876 59276
rect 426979 32240 433851 39173
rect 306753 26209 313014 27651
<< metal5 >>
rect 166394 703100 171394 704800
rect 176694 703100 181694 704800
rect 218094 703100 223094 704800
rect 228394 703100 233394 704800
rect 319794 703100 324794 704800
rect 330094 703100 335094 704800
rect 516238 698932 521238 699090
rect 516238 696670 516456 698932
rect 515321 693856 516456 696670
rect 520966 696670 521238 698932
rect 520966 693856 522787 696670
rect 515321 672866 522787 693856
rect 106520 665257 280703 672722
rect 106520 561595 114019 665257
rect 6412 560186 114019 561595
rect 3942 560048 114019 560186
rect 3942 555362 4066 560048
rect 9170 555362 114019 560048
rect 3942 555186 114019 555362
rect 6412 554130 114019 555186
rect 106520 475380 114019 554130
rect 106520 470309 106611 475380
rect 113894 470309 114019 475380
rect 106520 455661 114019 470309
rect 106520 454319 106619 455661
rect 113903 454319 114019 455661
rect 106520 441575 114019 454319
rect 106520 440408 106630 441575
rect 113902 440408 114019 441575
rect 106520 313538 114019 440408
rect 106520 310456 106704 313538
rect 113848 310456 114019 313538
rect 106520 280018 114019 310456
rect 106520 278712 106628 280018
rect 113928 278712 114019 280018
rect 106520 232157 114019 278712
rect 106520 224846 106878 232157
rect 113676 224846 114019 232157
rect 106520 224434 114019 224846
rect 150783 571845 169318 579095
rect 150783 489095 158033 571845
rect 150783 481845 169318 489095
rect 150783 462824 158033 481845
rect 150783 461395 150899 462824
rect 157916 461395 158033 462824
rect 150783 440395 158033 461395
rect 150783 439040 150941 440395
rect 157881 439040 158033 440395
rect 150783 399095 158033 439040
rect 150783 391845 169318 399095
rect 150783 309095 158033 391845
rect 150783 301845 169318 309095
rect 150783 219095 158033 301845
rect 150783 216733 169318 219095
rect 8595 215634 169318 216733
rect 4098 215436 169318 215634
rect 4098 210800 4232 215436
rect 9414 211845 169318 215436
rect 9414 210800 158033 211845
rect 4098 210634 158033 210800
rect 8595 209483 158033 210634
rect 106520 201306 114019 201663
rect 106520 194909 106922 201306
rect 113632 194909 114019 201306
rect 106520 139242 114019 194909
rect 106520 138416 106578 139242
rect 113928 138416 114019 139242
rect 106520 59276 114019 138416
rect 106520 58454 106648 59276
rect 113876 58454 114019 59276
rect 106520 18754 114019 58454
rect 150783 129095 158033 209483
rect 150783 121845 169318 129095
rect 150783 39095 158033 121845
rect 150783 31845 169318 39095
rect 273238 31207 280703 665257
rect 305969 665400 522787 672866
rect 305969 281232 313435 665400
rect 418431 572089 434054 579339
rect 426804 546276 434054 572089
rect 466215 577278 473681 665400
rect 466215 569837 466468 577278
rect 473449 569837 473681 577278
rect 466215 560021 473681 569837
rect 466215 553646 466599 560021
rect 473439 553646 473681 560021
rect 466215 553211 473681 553646
rect 553960 551280 577018 551988
rect 553960 550970 580932 551280
rect 553960 546532 575622 550970
rect 580746 546532 580932 550970
rect 553960 546280 580932 546532
rect 553960 546276 577018 546280
rect 426804 544738 577018 546276
rect 426804 539026 561210 544738
rect 426804 489339 434054 539026
rect 418431 482089 434054 489339
rect 426804 399339 434054 482089
rect 466215 530621 473681 530943
rect 466215 523885 466547 530621
rect 473413 523885 473681 530621
rect 466215 412769 473681 523885
rect 466206 412620 473703 412769
rect 466206 410038 466355 412620
rect 473541 410038 473703 412620
rect 466206 409865 473703 410038
rect 418431 392089 434054 399339
rect 426804 309339 434054 392089
rect 418431 302089 434054 309339
rect 426804 298253 434054 302089
rect 322531 298063 434054 298253
rect 322531 293627 322730 298063
rect 326798 293627 434054 298063
rect 322531 293461 434054 293627
rect 305969 279800 306274 281232
rect 312971 279800 313435 281232
rect 305969 27651 313435 279800
rect 426804 237151 434054 293461
rect 466215 255107 473681 409865
rect 466215 247031 466498 255107
rect 473424 247031 473681 255107
rect 466215 246663 473681 247031
rect 426804 235850 577018 237151
rect 426804 235522 580166 235850
rect 426804 231084 574962 235522
rect 580086 231084 580166 235522
rect 426804 230850 580166 231084
rect 426804 229901 577018 230850
rect 426804 219339 434054 229901
rect 418431 212089 434054 219339
rect 426804 129339 434054 212089
rect 418431 122089 434054 129339
rect 426804 39339 434054 122089
rect 418431 39173 434054 39339
rect 418431 32240 426979 39173
rect 433851 32240 434054 39173
rect 418431 32089 434054 32240
rect 466215 221314 473681 221672
rect 466215 211313 466529 221314
rect 473424 211313 473681 221314
rect 466215 149329 473681 211313
rect 466215 147502 578773 149329
rect 466215 147254 580654 147502
rect 466215 142816 575132 147254
rect 580256 142816 580654 147254
rect 466215 142502 580654 142816
rect 466215 141863 578773 142502
rect 305969 26209 306753 27651
rect 313014 26209 313435 27651
rect 305969 26129 313435 26209
rect 466215 26129 473681 141863
rect 305969 18663 473687 26129
<< comment >>
rect 0 704800 585600 705600
rect 0 800 800 704800
rect 533438 596264 551793 600607
rect 27798 503403 49688 511786
rect 18736 437627 38275 444818
rect 533336 425671 556320 432270
rect 533020 363414 550674 368496
rect 560302 365830 579683 368729
rect 55678 334437 70405 337219
rect 513224 325832 535292 331582
rect 16454 272114 23660 275184
rect 15452 135036 29200 138506
rect 518574 124676 539974 129892
rect 11782 61490 26398 65162
rect 584800 800 585600 704800
rect 0 0 585600 800
use analog_mux_sel1v8  analog_mux_sel1v8_0
timestamp 1713903757
transform 0 -1 583347 1 0 361407
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_1
timestamp 1713903757
transform 0 1 5348 1 0 462156
box -5530 -288 4452 6736
use analog_mux_sel1v8  analog_mux_sel1v8_2
timestamp 1713903757
transform -1 0 6199 0 1 427752
box -5530 -288 4452 6736
use bias_generator  bias_generator_0
timestamp 1713896310
transform 0 -1 291742 1 0 33373
box -902 -6353 245156 3114
use lpopamp  lpopamp_0 ../../chipalooza/sky130_rodovalho_ip__lpopamp/mag
timestamp 1713038477
transform 0 1 537526 1 0 246598
box -7000 0 81800 36300
use power_stage  power_stage_0
array 0 6 90000 0 0 -111006
timestamp 1713809566
transform 0 -1 234941 1 0 120408
box -89200 -44204 -9499 66802
use power_stage  power_stage_1
array 0 6 90000 0 0 111006
timestamp 1713809566
transform 0 1 351850 1 0 120408
box -89200 -44204 -9499 66802
use SDC  SDC_0
timestamp 1541985909
transform 1 0 536101 0 1 95480
box -29735 -18309 17962 24495
use sky130_ajc_ip__brownout  sky130_ajc_ip__brownout_0 ../../chipalooza/sky130_ajc_ip__brownout/mag
timestamp 1713419710
transform 0 1 33740 -1 0 89134
box -1604 -1987 43293 41283
use sky130_ajc_ip__overvoltage  sky130_ajc_ip__overvoltage_0 ../../chipalooza/sky130_ajc_ip__overvoltage/mag
timestamp 1713210720
transform 0 1 34176 -1 0 156926
box -2433 -2390 42464 28880
use sky130_ajc_ip__por  sky130_ajc_ip__por_0 ../../chipalooza/sky130_ajc_ip__por/mag
timestamp 1713454396
transform 0 1 28804 -1 0 294712
box -1604 -1987 43293 41283
use sky130_ak_ip__comparator  sky130_ak_ip__comparator_0 ../../chipalooza/sky130_ak_ip__comparator/mag
timestamp 1713602081
transform 0 -1 18376 1 0 319360
box -1900 -33700 39700 13700
use sky130_be_ip__lsxo  sky130_be_ip__lsxo_0 ../../chipalooza/sky130_be_ip__lsxo/mag
timestamp 1713362978
transform 0 -1 558491 1 0 410746
box 1626 -23704 25570 -812
use sky130_ht_ip__hsxo_cpz1  sky130_ht_ip__hsxo_cpz1_0 ../../chipalooza/hsxo-cpz1/mag
timestamp 1713816941
transform -1 0 569204 0 1 342778
box -3162 -7320 32492 17749
use sky130_od_ip__tempsensor_ext_vp  sky130_od_ip__tempsensor_ext_vp_0 ../../chipalooza/sky130_od_ip__tempsensor/mag
timestamp 1713856378
transform 1 0 9095 0 1 442073
box -584 -5030 6610 3202
use sky130_td_ip__opamp_hp  sky130_td_ip__opamp_hp_0 ../../chipalooza/sky130_td_ip__opamp_hp/mag
timestamp 1713675868
transform 0 1 10847 1 0 489761
box -7724 -6929 51340 16206
use sky130_vbl_ip__overvoltage  sky130_vbl_ip__overvoltage_0 ../../chipalooza/sky130_vbl_ip__overvoltage/mag
timestamp 1713724750
transform 1 0 539503 0 1 576713
box -18218 -4002 24405 17489
<< labels >>
flabel metal3 s 800 681042 2500 686042 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 800 644642 2460 649442 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 800 634642 2460 639442 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 800 205688 2460 210488 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 800 215688 2460 220488 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 800 560242 2460 565042 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 800 550242 2460 555042 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 800 173688 2460 178488 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 800 163688 2460 168488 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal4 15162 171077 15162 171077 0 FreeSans 16000 0 0 0 vssd2
flabel metal4 13496 642110 13496 642110 0 FreeSans 16000 0 0 0 vccd2
flabel comment 542585 598389 542585 598389 0 FreeSans 16000 0 0 0 overvoltage
flabel comment 544548 428758 544548 428758 0 FreeSans 16000 0 0 0 LSXO
flabel metal4 26979 17673 26979 17673 0 FreeSans 16000 0 0 0 bias_reference_voltage
flabel comment 569786 367507 569796 367507 0 FreeSans 16000 0 0 0 1.2V_reference
flabel comment 29461 503602 46827 511520 0 FreeSans 16000 0 0 0 HGBW_op_amp
flabel comment 29455 441019 29455 441019 0 FreeSans 16000 0 0 0 temp_sensor
flabel comment 63088 335906 63088 335906 0 FreeSans 16000 0 0 0 comparator
flabel comment 19790 273514 19790 273514 0 FreeSans 16000 0 0 0 por
flabel comment 22326 136704 22326 136704 0 FreeSans 16000 0 0 0 overvoltage
flabel comment 18856 63292 18856 63292 0 FreeSans 16000 0 0 0 brownout
flabel comment 530076 127352 530076 127352 0 FreeSans 16000 0 0 0 temp_sensor
flabel comment 541846 366090 541846 366090 0 FreeSans 16000 0 0 0 HSXO
flabel comment 524460 328506 524460 328506 0 FreeSans 16000 0 0 0 LP_op_amp
<< end >>
